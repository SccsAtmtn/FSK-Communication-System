module rHammingCode(datain, dataout);

wire [7:0] hamming[4095:0];
assign hamming[0] = 8'b00000000;
assign hamming[1] = 8'b00000000;
assign hamming[2] = 8'b00000000;
assign hamming[3] = 8'b00000001;
assign hamming[4] = 8'b00000000;
assign hamming[5] = 8'b00000001;
assign hamming[6] = 8'b00000001;
assign hamming[7] = 8'b00000001;
assign hamming[8] = 8'b00000000;
assign hamming[9] = 8'b00000010;
assign hamming[10] = 8'b00000100;
assign hamming[11] = 8'b00001000;
assign hamming[12] = 8'b00001001;
assign hamming[13] = 8'b00000101;
assign hamming[14] = 8'b00000011;
assign hamming[15] = 8'b00000001;
assign hamming[16] = 8'b00000000;
assign hamming[17] = 8'b00000010;
assign hamming[18] = 8'b00001010;
assign hamming[19] = 8'b00000110;
assign hamming[20] = 8'b00000111;
assign hamming[21] = 8'b00001011;
assign hamming[22] = 8'b00000011;
assign hamming[23] = 8'b00000001;
assign hamming[24] = 8'b00000010;
assign hamming[25] = 8'b00000010;
assign hamming[26] = 8'b00000011;
assign hamming[27] = 8'b00000010;
assign hamming[28] = 8'b00000011;
assign hamming[29] = 8'b00000010;
assign hamming[30] = 8'b00000011;
assign hamming[31] = 8'b00000011;
assign hamming[32] = 8'b00000000;
assign hamming[33] = 8'b00001100;
assign hamming[34] = 8'b00000100;
assign hamming[35] = 8'b00000110;
assign hamming[36] = 8'b00000111;
assign hamming[37] = 8'b00000101;
assign hamming[38] = 8'b00001101;
assign hamming[39] = 8'b00000001;
assign hamming[40] = 8'b00000100;
assign hamming[41] = 8'b00000101;
assign hamming[42] = 8'b00000100;
assign hamming[43] = 8'b00000100;
assign hamming[44] = 8'b00000101;
assign hamming[45] = 8'b00000101;
assign hamming[46] = 8'b00000100;
assign hamming[47] = 8'b00000101;
assign hamming[48] = 8'b00000111;
assign hamming[49] = 8'b00000110;
assign hamming[50] = 8'b00000110;
assign hamming[51] = 8'b00000110;
assign hamming[52] = 8'b00000111;
assign hamming[53] = 8'b00000111;
assign hamming[54] = 8'b00000111;
assign hamming[55] = 8'b00000110;
assign hamming[56] = 8'b00001110;
assign hamming[57] = 8'b00000010;
assign hamming[58] = 8'b00000100;
assign hamming[59] = 8'b00000110;
assign hamming[60] = 8'b00000111;
assign hamming[61] = 8'b00000101;
assign hamming[62] = 8'b00000011;
assign hamming[63] = 8'b00001111;
assign hamming[64] = 8'b00000000;
assign hamming[65] = 8'b00001100;
assign hamming[66] = 8'b00001010;
assign hamming[67] = 8'b00001000;
assign hamming[68] = 8'b00001001;
assign hamming[69] = 8'b00001011;
assign hamming[70] = 8'b00001101;
assign hamming[71] = 8'b00000001;
assign hamming[72] = 8'b00001001;
assign hamming[73] = 8'b00001000;
assign hamming[74] = 8'b00001000;
assign hamming[75] = 8'b00001000;
assign hamming[76] = 8'b00001001;
assign hamming[77] = 8'b00001001;
assign hamming[78] = 8'b00001001;
assign hamming[79] = 8'b00001000;
assign hamming[80] = 8'b00001010;
assign hamming[81] = 8'b00001011;
assign hamming[82] = 8'b00001010;
assign hamming[83] = 8'b00001010;
assign hamming[84] = 8'b00001011;
assign hamming[85] = 8'b00001011;
assign hamming[86] = 8'b00001010;
assign hamming[87] = 8'b00001011;
assign hamming[88] = 8'b00001110;
assign hamming[89] = 8'b00000010;
assign hamming[90] = 8'b00001010;
assign hamming[91] = 8'b00001000;
assign hamming[92] = 8'b00001001;
assign hamming[93] = 8'b00001011;
assign hamming[94] = 8'b00000011;
assign hamming[95] = 8'b00001111;
assign hamming[96] = 8'b00001100;
assign hamming[97] = 8'b00001100;
assign hamming[98] = 8'b00001101;
assign hamming[99] = 8'b00001100;
assign hamming[100] = 8'b00001101;
assign hamming[101] = 8'b00001100;
assign hamming[102] = 8'b00001101;
assign hamming[103] = 8'b00001101;
assign hamming[104] = 8'b00001110;
assign hamming[105] = 8'b00001100;
assign hamming[106] = 8'b00000100;
assign hamming[107] = 8'b00001000;
assign hamming[108] = 8'b00001001;
assign hamming[109] = 8'b00000101;
assign hamming[110] = 8'b00001101;
assign hamming[111] = 8'b00001111;
assign hamming[112] = 8'b00001110;
assign hamming[113] = 8'b00001100;
assign hamming[114] = 8'b00001010;
assign hamming[115] = 8'b00000110;
assign hamming[116] = 8'b00000111;
assign hamming[117] = 8'b00001011;
assign hamming[118] = 8'b00001101;
assign hamming[119] = 8'b00001111;
assign hamming[120] = 8'b00001110;
assign hamming[121] = 8'b00001110;
assign hamming[122] = 8'b00001110;
assign hamming[123] = 8'b00001111;
assign hamming[124] = 8'b00001110;
assign hamming[125] = 8'b00001111;
assign hamming[126] = 8'b00001111;
assign hamming[127] = 8'b00001111;
assign hamming[128] = 8'b00000000;
assign hamming[129] = 8'b00010000;
assign hamming[130] = 8'b00100000;
assign hamming[131] = 8'b01000000;
assign hamming[132] = 8'b01000001;
assign hamming[133] = 8'b00100001;
assign hamming[134] = 8'b00010001;
assign hamming[135] = 8'b00000001;
assign hamming[136] = 8'b10000000;
assign hamming[137] = 8'b11111111;
assign hamming[138] = 8'b11111111;
assign hamming[139] = 8'b11111111;
assign hamming[140] = 8'b11111111;
assign hamming[141] = 8'b11111111;
assign hamming[142] = 8'b11111111;
assign hamming[143] = 8'b10000001;
assign hamming[144] = 8'b11111111;
assign hamming[145] = 8'b10000010;
assign hamming[146] = 8'b11111111;
assign hamming[147] = 8'b11111111;
assign hamming[148] = 8'b11111111;
assign hamming[149] = 8'b11111111;
assign hamming[150] = 8'b10000011;
assign hamming[151] = 8'b11111111;
assign hamming[152] = 8'b00010010;
assign hamming[153] = 8'b00000010;
assign hamming[154] = 8'b01000010;
assign hamming[155] = 8'b00100010;
assign hamming[156] = 8'b00100011;
assign hamming[157] = 8'b01000011;
assign hamming[158] = 8'b00000011;
assign hamming[159] = 8'b00010011;
assign hamming[160] = 8'b11111111;
assign hamming[161] = 8'b11111111;
assign hamming[162] = 8'b10000100;
assign hamming[163] = 8'b11111111;
assign hamming[164] = 8'b11111111;
assign hamming[165] = 8'b10000101;
assign hamming[166] = 8'b11111111;
assign hamming[167] = 8'b11111111;
assign hamming[168] = 8'b00100100;
assign hamming[169] = 8'b01000100;
assign hamming[170] = 8'b00000100;
assign hamming[171] = 8'b00010100;
assign hamming[172] = 8'b00010101;
assign hamming[173] = 8'b00000101;
assign hamming[174] = 8'b01000101;
assign hamming[175] = 8'b00100101;
assign hamming[176] = 8'b01000110;
assign hamming[177] = 8'b00100110;
assign hamming[178] = 8'b00010110;
assign hamming[179] = 8'b00000110;
assign hamming[180] = 8'b00000111;
assign hamming[181] = 8'b00010111;
assign hamming[182] = 8'b00100111;
assign hamming[183] = 8'b01000111;
assign hamming[184] = 8'b11111111;
assign hamming[185] = 8'b11111111;
assign hamming[186] = 8'b11111111;
assign hamming[187] = 8'b10000110;
assign hamming[188] = 8'b10000111;
assign hamming[189] = 8'b11111111;
assign hamming[190] = 8'b11111111;
assign hamming[191] = 8'b11111111;
assign hamming[192] = 8'b11111111;
assign hamming[193] = 8'b11111111;
assign hamming[194] = 8'b11111111;
assign hamming[195] = 8'b10001000;
assign hamming[196] = 8'b10001001;
assign hamming[197] = 8'b11111111;
assign hamming[198] = 8'b11111111;
assign hamming[199] = 8'b11111111;
assign hamming[200] = 8'b01001000;
assign hamming[201] = 8'b00101000;
assign hamming[202] = 8'b00011000;
assign hamming[203] = 8'b00001000;
assign hamming[204] = 8'b00001001;
assign hamming[205] = 8'b00011001;
assign hamming[206] = 8'b00101001;
assign hamming[207] = 8'b01001001;
assign hamming[208] = 8'b00101010;
assign hamming[209] = 8'b01001010;
assign hamming[210] = 8'b00001010;
assign hamming[211] = 8'b00011010;
assign hamming[212] = 8'b00011011;
assign hamming[213] = 8'b00001011;
assign hamming[214] = 8'b01001011;
assign hamming[215] = 8'b00101011;
assign hamming[216] = 8'b11111111;
assign hamming[217] = 8'b11111111;
assign hamming[218] = 8'b10001010;
assign hamming[219] = 8'b11111111;
assign hamming[220] = 8'b11111111;
assign hamming[221] = 8'b10001011;
assign hamming[222] = 8'b11111111;
assign hamming[223] = 8'b11111111;
assign hamming[224] = 8'b00011100;
assign hamming[225] = 8'b00001100;
assign hamming[226] = 8'b01001100;
assign hamming[227] = 8'b00101100;
assign hamming[228] = 8'b00101101;
assign hamming[229] = 8'b01001101;
assign hamming[230] = 8'b00001101;
assign hamming[231] = 8'b00011101;
assign hamming[232] = 8'b11111111;
assign hamming[233] = 8'b10001100;
assign hamming[234] = 8'b11111111;
assign hamming[235] = 8'b11111111;
assign hamming[236] = 8'b11111111;
assign hamming[237] = 8'b11111111;
assign hamming[238] = 8'b10001101;
assign hamming[239] = 8'b11111111;
assign hamming[240] = 8'b10001110;
assign hamming[241] = 8'b11111111;
assign hamming[242] = 8'b11111111;
assign hamming[243] = 8'b11111111;
assign hamming[244] = 8'b11111111;
assign hamming[245] = 8'b11111111;
assign hamming[246] = 8'b11111111;
assign hamming[247] = 8'b10001111;
assign hamming[248] = 8'b00001110;
assign hamming[249] = 8'b00011110;
assign hamming[250] = 8'b00101110;
assign hamming[251] = 8'b01001110;
assign hamming[252] = 8'b01001111;
assign hamming[253] = 8'b00101111;
assign hamming[254] = 8'b00011111;
assign hamming[255] = 8'b00001111;
assign hamming[256] = 8'b00000000;
assign hamming[257] = 8'b00010000;
assign hamming[258] = 8'b01010000;
assign hamming[259] = 8'b00110000;
assign hamming[260] = 8'b00110001;
assign hamming[261] = 8'b01010001;
assign hamming[262] = 8'b00010001;
assign hamming[263] = 8'b00000001;
assign hamming[264] = 8'b11111111;
assign hamming[265] = 8'b10010000;
assign hamming[266] = 8'b11111111;
assign hamming[267] = 8'b11111111;
assign hamming[268] = 8'b11111111;
assign hamming[269] = 8'b11111111;
assign hamming[270] = 8'b10010001;
assign hamming[271] = 8'b11111111;
assign hamming[272] = 8'b10010010;
assign hamming[273] = 8'b11111111;
assign hamming[274] = 8'b11111111;
assign hamming[275] = 8'b11111111;
assign hamming[276] = 8'b11111111;
assign hamming[277] = 8'b11111111;
assign hamming[278] = 8'b11111111;
assign hamming[279] = 8'b10010011;
assign hamming[280] = 8'b00010010;
assign hamming[281] = 8'b00000010;
assign hamming[282] = 8'b00110010;
assign hamming[283] = 8'b01010010;
assign hamming[284] = 8'b01010011;
assign hamming[285] = 8'b00110011;
assign hamming[286] = 8'b00000011;
assign hamming[287] = 8'b00010011;
assign hamming[288] = 8'b11111111;
assign hamming[289] = 8'b11111111;
assign hamming[290] = 8'b11111111;
assign hamming[291] = 8'b10010100;
assign hamming[292] = 8'b10010101;
assign hamming[293] = 8'b11111111;
assign hamming[294] = 8'b11111111;
assign hamming[295] = 8'b11111111;
assign hamming[296] = 8'b01010100;
assign hamming[297] = 8'b00110100;
assign hamming[298] = 8'b00000100;
assign hamming[299] = 8'b00010100;
assign hamming[300] = 8'b00010101;
assign hamming[301] = 8'b00000101;
assign hamming[302] = 8'b00110101;
assign hamming[303] = 8'b01010101;
assign hamming[304] = 8'b00110110;
assign hamming[305] = 8'b01010110;
assign hamming[306] = 8'b00010110;
assign hamming[307] = 8'b00000110;
assign hamming[308] = 8'b00000111;
assign hamming[309] = 8'b00010111;
assign hamming[310] = 8'b01010111;
assign hamming[311] = 8'b00110111;
assign hamming[312] = 8'b11111111;
assign hamming[313] = 8'b11111111;
assign hamming[314] = 8'b10010110;
assign hamming[315] = 8'b11111111;
assign hamming[316] = 8'b11111111;
assign hamming[317] = 8'b10010111;
assign hamming[318] = 8'b11111111;
assign hamming[319] = 8'b11111111;
assign hamming[320] = 8'b11111111;
assign hamming[321] = 8'b11111111;
assign hamming[322] = 8'b10011000;
assign hamming[323] = 8'b11111111;
assign hamming[324] = 8'b11111111;
assign hamming[325] = 8'b10011001;
assign hamming[326] = 8'b11111111;
assign hamming[327] = 8'b11111111;
assign hamming[328] = 8'b00111000;
assign hamming[329] = 8'b01011000;
assign hamming[330] = 8'b00011000;
assign hamming[331] = 8'b00001000;
assign hamming[332] = 8'b00001001;
assign hamming[333] = 8'b00011001;
assign hamming[334] = 8'b01011001;
assign hamming[335] = 8'b00111001;
assign hamming[336] = 8'b01011010;
assign hamming[337] = 8'b00111010;
assign hamming[338] = 8'b00001010;
assign hamming[339] = 8'b00011010;
assign hamming[340] = 8'b00011011;
assign hamming[341] = 8'b00001011;
assign hamming[342] = 8'b00111011;
assign hamming[343] = 8'b01011011;
assign hamming[344] = 8'b11111111;
assign hamming[345] = 8'b11111111;
assign hamming[346] = 8'b11111111;
assign hamming[347] = 8'b10011010;
assign hamming[348] = 8'b10011011;
assign hamming[349] = 8'b11111111;
assign hamming[350] = 8'b11111111;
assign hamming[351] = 8'b11111111;
assign hamming[352] = 8'b00011100;
assign hamming[353] = 8'b00001100;
assign hamming[354] = 8'b00111100;
assign hamming[355] = 8'b01011100;
assign hamming[356] = 8'b01011101;
assign hamming[357] = 8'b00111101;
assign hamming[358] = 8'b00001101;
assign hamming[359] = 8'b00011101;
assign hamming[360] = 8'b10011100;
assign hamming[361] = 8'b11111111;
assign hamming[362] = 8'b11111111;
assign hamming[363] = 8'b11111111;
assign hamming[364] = 8'b11111111;
assign hamming[365] = 8'b11111111;
assign hamming[366] = 8'b11111111;
assign hamming[367] = 8'b10011101;
assign hamming[368] = 8'b11111111;
assign hamming[369] = 8'b10011110;
assign hamming[370] = 8'b11111111;
assign hamming[371] = 8'b11111111;
assign hamming[372] = 8'b11111111;
assign hamming[373] = 8'b11111111;
assign hamming[374] = 8'b10011111;
assign hamming[375] = 8'b11111111;
assign hamming[376] = 8'b00001110;
assign hamming[377] = 8'b00011110;
assign hamming[378] = 8'b01011110;
assign hamming[379] = 8'b00111110;
assign hamming[380] = 8'b00111111;
assign hamming[381] = 8'b01011111;
assign hamming[382] = 8'b00011111;
assign hamming[383] = 8'b00001111;
assign hamming[384] = 8'b00010000;
assign hamming[385] = 8'b00010000;
assign hamming[386] = 8'b00010001;
assign hamming[387] = 8'b00010000;
assign hamming[388] = 8'b00010001;
assign hamming[389] = 8'b00010000;
assign hamming[390] = 8'b00010001;
assign hamming[391] = 8'b00010001;
assign hamming[392] = 8'b00010010;
assign hamming[393] = 8'b00010000;
assign hamming[394] = 8'b00011000;
assign hamming[395] = 8'b00010100;
assign hamming[396] = 8'b00010101;
assign hamming[397] = 8'b00011001;
assign hamming[398] = 8'b00010001;
assign hamming[399] = 8'b00010011;
assign hamming[400] = 8'b00010010;
assign hamming[401] = 8'b00010000;
assign hamming[402] = 8'b00010110;
assign hamming[403] = 8'b00011010;
assign hamming[404] = 8'b00011011;
assign hamming[405] = 8'b00010111;
assign hamming[406] = 8'b00010001;
assign hamming[407] = 8'b00010011;
assign hamming[408] = 8'b00010010;
assign hamming[409] = 8'b00010010;
assign hamming[410] = 8'b00010010;
assign hamming[411] = 8'b00010011;
assign hamming[412] = 8'b00010010;
assign hamming[413] = 8'b00010011;
assign hamming[414] = 8'b00010011;
assign hamming[415] = 8'b00010011;
assign hamming[416] = 8'b00011100;
assign hamming[417] = 8'b00010000;
assign hamming[418] = 8'b00010110;
assign hamming[419] = 8'b00010100;
assign hamming[420] = 8'b00010101;
assign hamming[421] = 8'b00010111;
assign hamming[422] = 8'b00010001;
assign hamming[423] = 8'b00011101;
assign hamming[424] = 8'b00010101;
assign hamming[425] = 8'b00010100;
assign hamming[426] = 8'b00010100;
assign hamming[427] = 8'b00010100;
assign hamming[428] = 8'b00010101;
assign hamming[429] = 8'b00010101;
assign hamming[430] = 8'b00010101;
assign hamming[431] = 8'b00010100;
assign hamming[432] = 8'b00010110;
assign hamming[433] = 8'b00010111;
assign hamming[434] = 8'b00010110;
assign hamming[435] = 8'b00010110;
assign hamming[436] = 8'b00010111;
assign hamming[437] = 8'b00010111;
assign hamming[438] = 8'b00010110;
assign hamming[439] = 8'b00010111;
assign hamming[440] = 8'b00010010;
assign hamming[441] = 8'b00011110;
assign hamming[442] = 8'b00010110;
assign hamming[443] = 8'b00010100;
assign hamming[444] = 8'b00010101;
assign hamming[445] = 8'b00010111;
assign hamming[446] = 8'b00011111;
assign hamming[447] = 8'b00010011;
assign hamming[448] = 8'b00011100;
assign hamming[449] = 8'b00010000;
assign hamming[450] = 8'b00011000;
assign hamming[451] = 8'b00011010;
assign hamming[452] = 8'b00011011;
assign hamming[453] = 8'b00011001;
assign hamming[454] = 8'b00010001;
assign hamming[455] = 8'b00011101;
assign hamming[456] = 8'b00011000;
assign hamming[457] = 8'b00011001;
assign hamming[458] = 8'b00011000;
assign hamming[459] = 8'b00011000;
assign hamming[460] = 8'b00011001;
assign hamming[461] = 8'b00011001;
assign hamming[462] = 8'b00011000;
assign hamming[463] = 8'b00011001;
assign hamming[464] = 8'b00011011;
assign hamming[465] = 8'b00011010;
assign hamming[466] = 8'b00011010;
assign hamming[467] = 8'b00011010;
assign hamming[468] = 8'b00011011;
assign hamming[469] = 8'b00011011;
assign hamming[470] = 8'b00011011;
assign hamming[471] = 8'b00011010;
assign hamming[472] = 8'b00010010;
assign hamming[473] = 8'b00011110;
assign hamming[474] = 8'b00011000;
assign hamming[475] = 8'b00011010;
assign hamming[476] = 8'b00011011;
assign hamming[477] = 8'b00011001;
assign hamming[478] = 8'b00011111;
assign hamming[479] = 8'b00010011;
assign hamming[480] = 8'b00011100;
assign hamming[481] = 8'b00011100;
assign hamming[482] = 8'b00011100;
assign hamming[483] = 8'b00011101;
assign hamming[484] = 8'b00011100;
assign hamming[485] = 8'b00011101;
assign hamming[486] = 8'b00011101;
assign hamming[487] = 8'b00011101;
assign hamming[488] = 8'b00011100;
assign hamming[489] = 8'b00011110;
assign hamming[490] = 8'b00011000;
assign hamming[491] = 8'b00010100;
assign hamming[492] = 8'b00010101;
assign hamming[493] = 8'b00011001;
assign hamming[494] = 8'b00011111;
assign hamming[495] = 8'b00011101;
assign hamming[496] = 8'b00011100;
assign hamming[497] = 8'b00011110;
assign hamming[498] = 8'b00010110;
assign hamming[499] = 8'b00011010;
assign hamming[500] = 8'b00011011;
assign hamming[501] = 8'b00010111;
assign hamming[502] = 8'b00011111;
assign hamming[503] = 8'b00011101;
assign hamming[504] = 8'b00011110;
assign hamming[505] = 8'b00011110;
assign hamming[506] = 8'b00011111;
assign hamming[507] = 8'b00011110;
assign hamming[508] = 8'b00011111;
assign hamming[509] = 8'b00011110;
assign hamming[510] = 8'b00011111;
assign hamming[511] = 8'b00011111;
assign hamming[512] = 8'b00000000;
assign hamming[513] = 8'b01100000;
assign hamming[514] = 8'b00100000;
assign hamming[515] = 8'b00110000;
assign hamming[516] = 8'b00110001;
assign hamming[517] = 8'b00100001;
assign hamming[518] = 8'b01100001;
assign hamming[519] = 8'b00000001;
assign hamming[520] = 8'b11111111;
assign hamming[521] = 8'b11111111;
assign hamming[522] = 8'b10100000;
assign hamming[523] = 8'b11111111;
assign hamming[524] = 8'b11111111;
assign hamming[525] = 8'b10100001;
assign hamming[526] = 8'b11111111;
assign hamming[527] = 8'b11111111;
assign hamming[528] = 8'b11111111;
assign hamming[529] = 8'b11111111;
assign hamming[530] = 8'b11111111;
assign hamming[531] = 8'b10100010;
assign hamming[532] = 8'b10100011;
assign hamming[533] = 8'b11111111;
assign hamming[534] = 8'b11111111;
assign hamming[535] = 8'b11111111;
assign hamming[536] = 8'b01100010;
assign hamming[537] = 8'b00000010;
assign hamming[538] = 8'b00110010;
assign hamming[539] = 8'b00100010;
assign hamming[540] = 8'b00100011;
assign hamming[541] = 8'b00110011;
assign hamming[542] = 8'b00000011;
assign hamming[543] = 8'b01100011;
assign hamming[544] = 8'b10100100;
assign hamming[545] = 8'b11111111;
assign hamming[546] = 8'b11111111;
assign hamming[547] = 8'b11111111;
assign hamming[548] = 8'b11111111;
assign hamming[549] = 8'b11111111;
assign hamming[550] = 8'b11111111;
assign hamming[551] = 8'b10100101;
assign hamming[552] = 8'b00100100;
assign hamming[553] = 8'b00110100;
assign hamming[554] = 8'b00000100;
assign hamming[555] = 8'b01100100;
assign hamming[556] = 8'b01100101;
assign hamming[557] = 8'b00000101;
assign hamming[558] = 8'b00110101;
assign hamming[559] = 8'b00100101;
assign hamming[560] = 8'b00110110;
assign hamming[561] = 8'b00100110;
assign hamming[562] = 8'b01100110;
assign hamming[563] = 8'b00000110;
assign hamming[564] = 8'b00000111;
assign hamming[565] = 8'b01100111;
assign hamming[566] = 8'b00100111;
assign hamming[567] = 8'b00110111;
assign hamming[568] = 8'b11111111;
assign hamming[569] = 8'b10100110;
assign hamming[570] = 8'b11111111;
assign hamming[571] = 8'b11111111;
assign hamming[572] = 8'b11111111;
assign hamming[573] = 8'b11111111;
assign hamming[574] = 8'b10100111;
assign hamming[575] = 8'b11111111;
assign hamming[576] = 8'b11111111;
assign hamming[577] = 8'b10101000;
assign hamming[578] = 8'b11111111;
assign hamming[579] = 8'b11111111;
assign hamming[580] = 8'b11111111;
assign hamming[581] = 8'b11111111;
assign hamming[582] = 8'b10101001;
assign hamming[583] = 8'b11111111;
assign hamming[584] = 8'b00111000;
assign hamming[585] = 8'b00101000;
assign hamming[586] = 8'b01101000;
assign hamming[587] = 8'b00001000;
assign hamming[588] = 8'b00001001;
assign hamming[589] = 8'b01101001;
assign hamming[590] = 8'b00101001;
assign hamming[591] = 8'b00111001;
assign hamming[592] = 8'b00101010;
assign hamming[593] = 8'b00111010;
assign hamming[594] = 8'b00001010;
assign hamming[595] = 8'b01101010;
assign hamming[596] = 8'b01101011;
assign hamming[597] = 8'b00001011;
assign hamming[598] = 8'b00111011;
assign hamming[599] = 8'b00101011;
assign hamming[600] = 8'b10101010;
assign hamming[601] = 8'b11111111;
assign hamming[602] = 8'b11111111;
assign hamming[603] = 8'b11111111;
assign hamming[604] = 8'b11111111;
assign hamming[605] = 8'b11111111;
assign hamming[606] = 8'b11111111;
assign hamming[607] = 8'b10101011;
assign hamming[608] = 8'b01101100;
assign hamming[609] = 8'b00001100;
assign hamming[610] = 8'b00111100;
assign hamming[611] = 8'b00101100;
assign hamming[612] = 8'b00101101;
assign hamming[613] = 8'b00111101;
assign hamming[614] = 8'b00001101;
assign hamming[615] = 8'b01101101;
assign hamming[616] = 8'b11111111;
assign hamming[617] = 8'b11111111;
assign hamming[618] = 8'b11111111;
assign hamming[619] = 8'b10101100;
assign hamming[620] = 8'b10101101;
assign hamming[621] = 8'b11111111;
assign hamming[622] = 8'b11111111;
assign hamming[623] = 8'b11111111;
assign hamming[624] = 8'b11111111;
assign hamming[625] = 8'b11111111;
assign hamming[626] = 8'b10101110;
assign hamming[627] = 8'b11111111;
assign hamming[628] = 8'b11111111;
assign hamming[629] = 8'b10101111;
assign hamming[630] = 8'b11111111;
assign hamming[631] = 8'b11111111;
assign hamming[632] = 8'b00001110;
assign hamming[633] = 8'b01101110;
assign hamming[634] = 8'b00101110;
assign hamming[635] = 8'b00111110;
assign hamming[636] = 8'b00111111;
assign hamming[637] = 8'b00101111;
assign hamming[638] = 8'b01101111;
assign hamming[639] = 8'b00001111;
assign hamming[640] = 8'b00100000;
assign hamming[641] = 8'b00100001;
assign hamming[642] = 8'b00100000;
assign hamming[643] = 8'b00100000;
assign hamming[644] = 8'b00100001;
assign hamming[645] = 8'b00100001;
assign hamming[646] = 8'b00100000;
assign hamming[647] = 8'b00100001;
assign hamming[648] = 8'b00100100;
assign hamming[649] = 8'b00101000;
assign hamming[650] = 8'b00100000;
assign hamming[651] = 8'b00100010;
assign hamming[652] = 8'b00100011;
assign hamming[653] = 8'b00100001;
assign hamming[654] = 8'b00101001;
assign hamming[655] = 8'b00100101;
assign hamming[656] = 8'b00101010;
assign hamming[657] = 8'b00100110;
assign hamming[658] = 8'b00100000;
assign hamming[659] = 8'b00100010;
assign hamming[660] = 8'b00100011;
assign hamming[661] = 8'b00100001;
assign hamming[662] = 8'b00100111;
assign hamming[663] = 8'b00101011;
assign hamming[664] = 8'b00100011;
assign hamming[665] = 8'b00100010;
assign hamming[666] = 8'b00100010;
assign hamming[667] = 8'b00100010;
assign hamming[668] = 8'b00100011;
assign hamming[669] = 8'b00100011;
assign hamming[670] = 8'b00100011;
assign hamming[671] = 8'b00100010;
assign hamming[672] = 8'b00100100;
assign hamming[673] = 8'b00100110;
assign hamming[674] = 8'b00100000;
assign hamming[675] = 8'b00101100;
assign hamming[676] = 8'b00101101;
assign hamming[677] = 8'b00100001;
assign hamming[678] = 8'b00100111;
assign hamming[679] = 8'b00100101;
assign hamming[680] = 8'b00100100;
assign hamming[681] = 8'b00100100;
assign hamming[682] = 8'b00100100;
assign hamming[683] = 8'b00100101;
assign hamming[684] = 8'b00100100;
assign hamming[685] = 8'b00100101;
assign hamming[686] = 8'b00100101;
assign hamming[687] = 8'b00100101;
assign hamming[688] = 8'b00100110;
assign hamming[689] = 8'b00100110;
assign hamming[690] = 8'b00100111;
assign hamming[691] = 8'b00100110;
assign hamming[692] = 8'b00100111;
assign hamming[693] = 8'b00100110;
assign hamming[694] = 8'b00100111;
assign hamming[695] = 8'b00100111;
assign hamming[696] = 8'b00100100;
assign hamming[697] = 8'b00100110;
assign hamming[698] = 8'b00101110;
assign hamming[699] = 8'b00100010;
assign hamming[700] = 8'b00100011;
assign hamming[701] = 8'b00101111;
assign hamming[702] = 8'b00100111;
assign hamming[703] = 8'b00100101;
assign hamming[704] = 8'b00101010;
assign hamming[705] = 8'b00101000;
assign hamming[706] = 8'b00100000;
assign hamming[707] = 8'b00101100;
assign hamming[708] = 8'b00101101;
assign hamming[709] = 8'b00100001;
assign hamming[710] = 8'b00101001;
assign hamming[711] = 8'b00101011;
assign hamming[712] = 8'b00101000;
assign hamming[713] = 8'b00101000;
assign hamming[714] = 8'b00101001;
assign hamming[715] = 8'b00101000;
assign hamming[716] = 8'b00101001;
assign hamming[717] = 8'b00101000;
assign hamming[718] = 8'b00101001;
assign hamming[719] = 8'b00101001;
assign hamming[720] = 8'b00101010;
assign hamming[721] = 8'b00101010;
assign hamming[722] = 8'b00101010;
assign hamming[723] = 8'b00101011;
assign hamming[724] = 8'b00101010;
assign hamming[725] = 8'b00101011;
assign hamming[726] = 8'b00101011;
assign hamming[727] = 8'b00101011;
assign hamming[728] = 8'b00101010;
assign hamming[729] = 8'b00101000;
assign hamming[730] = 8'b00101110;
assign hamming[731] = 8'b00100010;
assign hamming[732] = 8'b00100011;
assign hamming[733] = 8'b00101111;
assign hamming[734] = 8'b00101001;
assign hamming[735] = 8'b00101011;
assign hamming[736] = 8'b00101101;
assign hamming[737] = 8'b00101100;
assign hamming[738] = 8'b00101100;
assign hamming[739] = 8'b00101100;
assign hamming[740] = 8'b00101101;
assign hamming[741] = 8'b00101101;
assign hamming[742] = 8'b00101101;
assign hamming[743] = 8'b00101100;
assign hamming[744] = 8'b00100100;
assign hamming[745] = 8'b00101000;
assign hamming[746] = 8'b00101110;
assign hamming[747] = 8'b00101100;
assign hamming[748] = 8'b00101101;
assign hamming[749] = 8'b00101111;
assign hamming[750] = 8'b00101001;
assign hamming[751] = 8'b00100101;
assign hamming[752] = 8'b00101010;
assign hamming[753] = 8'b00100110;
assign hamming[754] = 8'b00101110;
assign hamming[755] = 8'b00101100;
assign hamming[756] = 8'b00101101;
assign hamming[757] = 8'b00101111;
assign hamming[758] = 8'b00100111;
assign hamming[759] = 8'b00101011;
assign hamming[760] = 8'b00101110;
assign hamming[761] = 8'b00101111;
assign hamming[762] = 8'b00101110;
assign hamming[763] = 8'b00101110;
assign hamming[764] = 8'b00101111;
assign hamming[765] = 8'b00101111;
assign hamming[766] = 8'b00101110;
assign hamming[767] = 8'b00101111;
assign hamming[768] = 8'b00110001;
assign hamming[769] = 8'b00110000;
assign hamming[770] = 8'b00110000;
assign hamming[771] = 8'b00110000;
assign hamming[772] = 8'b00110001;
assign hamming[773] = 8'b00110001;
assign hamming[774] = 8'b00110001;
assign hamming[775] = 8'b00110000;
assign hamming[776] = 8'b00111000;
assign hamming[777] = 8'b00110100;
assign hamming[778] = 8'b00110010;
assign hamming[779] = 8'b00110000;
assign hamming[780] = 8'b00110001;
assign hamming[781] = 8'b00110011;
assign hamming[782] = 8'b00110101;
assign hamming[783] = 8'b00111001;
assign hamming[784] = 8'b00110110;
assign hamming[785] = 8'b00111010;
assign hamming[786] = 8'b00110010;
assign hamming[787] = 8'b00110000;
assign hamming[788] = 8'b00110001;
assign hamming[789] = 8'b00110011;
assign hamming[790] = 8'b00111011;
assign hamming[791] = 8'b00110111;
assign hamming[792] = 8'b00110010;
assign hamming[793] = 8'b00110011;
assign hamming[794] = 8'b00110010;
assign hamming[795] = 8'b00110010;
assign hamming[796] = 8'b00110011;
assign hamming[797] = 8'b00110011;
assign hamming[798] = 8'b00110010;
assign hamming[799] = 8'b00110011;
assign hamming[800] = 8'b00110110;
assign hamming[801] = 8'b00110100;
assign hamming[802] = 8'b00111100;
assign hamming[803] = 8'b00110000;
assign hamming[804] = 8'b00110001;
assign hamming[805] = 8'b00111101;
assign hamming[806] = 8'b00110101;
assign hamming[807] = 8'b00110111;
assign hamming[808] = 8'b00110100;
assign hamming[809] = 8'b00110100;
assign hamming[810] = 8'b00110101;
assign hamming[811] = 8'b00110100;
assign hamming[812] = 8'b00110101;
assign hamming[813] = 8'b00110100;
assign hamming[814] = 8'b00110101;
assign hamming[815] = 8'b00110101;
assign hamming[816] = 8'b00110110;
assign hamming[817] = 8'b00110110;
assign hamming[818] = 8'b00110110;
assign hamming[819] = 8'b00110111;
assign hamming[820] = 8'b00110110;
assign hamming[821] = 8'b00110111;
assign hamming[822] = 8'b00110111;
assign hamming[823] = 8'b00110111;
assign hamming[824] = 8'b00110110;
assign hamming[825] = 8'b00110100;
assign hamming[826] = 8'b00110010;
assign hamming[827] = 8'b00111110;
assign hamming[828] = 8'b00111111;
assign hamming[829] = 8'b00110011;
assign hamming[830] = 8'b00110101;
assign hamming[831] = 8'b00110111;
assign hamming[832] = 8'b00111000;
assign hamming[833] = 8'b00111010;
assign hamming[834] = 8'b00111100;
assign hamming[835] = 8'b00110000;
assign hamming[836] = 8'b00110001;
assign hamming[837] = 8'b00111101;
assign hamming[838] = 8'b00111011;
assign hamming[839] = 8'b00111001;
assign hamming[840] = 8'b00111000;
assign hamming[841] = 8'b00111000;
assign hamming[842] = 8'b00111000;
assign hamming[843] = 8'b00111001;
assign hamming[844] = 8'b00111000;
assign hamming[845] = 8'b00111001;
assign hamming[846] = 8'b00111001;
assign hamming[847] = 8'b00111001;
assign hamming[848] = 8'b00111010;
assign hamming[849] = 8'b00111010;
assign hamming[850] = 8'b00111011;
assign hamming[851] = 8'b00111010;
assign hamming[852] = 8'b00111011;
assign hamming[853] = 8'b00111010;
assign hamming[854] = 8'b00111011;
assign hamming[855] = 8'b00111011;
assign hamming[856] = 8'b00111000;
assign hamming[857] = 8'b00111010;
assign hamming[858] = 8'b00110010;
assign hamming[859] = 8'b00111110;
assign hamming[860] = 8'b00111111;
assign hamming[861] = 8'b00110011;
assign hamming[862] = 8'b00111011;
assign hamming[863] = 8'b00111001;
assign hamming[864] = 8'b00111100;
assign hamming[865] = 8'b00111101;
assign hamming[866] = 8'b00111100;
assign hamming[867] = 8'b00111100;
assign hamming[868] = 8'b00111101;
assign hamming[869] = 8'b00111101;
assign hamming[870] = 8'b00111100;
assign hamming[871] = 8'b00111101;
assign hamming[872] = 8'b00111000;
assign hamming[873] = 8'b00110100;
assign hamming[874] = 8'b00111100;
assign hamming[875] = 8'b00111110;
assign hamming[876] = 8'b00111111;
assign hamming[877] = 8'b00111101;
assign hamming[878] = 8'b00110101;
assign hamming[879] = 8'b00111001;
assign hamming[880] = 8'b00110110;
assign hamming[881] = 8'b00111010;
assign hamming[882] = 8'b00111100;
assign hamming[883] = 8'b00111110;
assign hamming[884] = 8'b00111111;
assign hamming[885] = 8'b00111101;
assign hamming[886] = 8'b00111011;
assign hamming[887] = 8'b00110111;
assign hamming[888] = 8'b00111111;
assign hamming[889] = 8'b00111110;
assign hamming[890] = 8'b00111110;
assign hamming[891] = 8'b00111110;
assign hamming[892] = 8'b00111111;
assign hamming[893] = 8'b00111111;
assign hamming[894] = 8'b00111111;
assign hamming[895] = 8'b00111110;
assign hamming[896] = 8'b01110000;
assign hamming[897] = 8'b00010000;
assign hamming[898] = 8'b00100000;
assign hamming[899] = 8'b00110000;
assign hamming[900] = 8'b00110001;
assign hamming[901] = 8'b00100001;
assign hamming[902] = 8'b00010001;
assign hamming[903] = 8'b01110001;
assign hamming[904] = 8'b11111111;
assign hamming[905] = 8'b11111111;
assign hamming[906] = 8'b11111111;
assign hamming[907] = 8'b10110000;
assign hamming[908] = 8'b10110001;
assign hamming[909] = 8'b11111111;
assign hamming[910] = 8'b11111111;
assign hamming[911] = 8'b11111111;
assign hamming[912] = 8'b11111111;
assign hamming[913] = 8'b11111111;
assign hamming[914] = 8'b10110010;
assign hamming[915] = 8'b11111111;
assign hamming[916] = 8'b11111111;
assign hamming[917] = 8'b10110011;
assign hamming[918] = 8'b11111111;
assign hamming[919] = 8'b11111111;
assign hamming[920] = 8'b00010010;
assign hamming[921] = 8'b01110010;
assign hamming[922] = 8'b00110010;
assign hamming[923] = 8'b00100010;
assign hamming[924] = 8'b00100011;
assign hamming[925] = 8'b00110011;
assign hamming[926] = 8'b01110011;
assign hamming[927] = 8'b00010011;
assign hamming[928] = 8'b11111111;
assign hamming[929] = 8'b10110100;
assign hamming[930] = 8'b11111111;
assign hamming[931] = 8'b11111111;
assign hamming[932] = 8'b11111111;
assign hamming[933] = 8'b11111111;
assign hamming[934] = 8'b10110101;
assign hamming[935] = 8'b11111111;
assign hamming[936] = 8'b00100100;
assign hamming[937] = 8'b00110100;
assign hamming[938] = 8'b01110100;
assign hamming[939] = 8'b00010100;
assign hamming[940] = 8'b00010101;
assign hamming[941] = 8'b01110101;
assign hamming[942] = 8'b00110101;
assign hamming[943] = 8'b00100101;
assign hamming[944] = 8'b00110110;
assign hamming[945] = 8'b00100110;
assign hamming[946] = 8'b00010110;
assign hamming[947] = 8'b01110110;
assign hamming[948] = 8'b01110111;
assign hamming[949] = 8'b00010111;
assign hamming[950] = 8'b00100111;
assign hamming[951] = 8'b00110111;
assign hamming[952] = 8'b10110110;
assign hamming[953] = 8'b11111111;
assign hamming[954] = 8'b11111111;
assign hamming[955] = 8'b11111111;
assign hamming[956] = 8'b11111111;
assign hamming[957] = 8'b11111111;
assign hamming[958] = 8'b11111111;
assign hamming[959] = 8'b10110111;
assign hamming[960] = 8'b10111000;
assign hamming[961] = 8'b11111111;
assign hamming[962] = 8'b11111111;
assign hamming[963] = 8'b11111111;
assign hamming[964] = 8'b11111111;
assign hamming[965] = 8'b11111111;
assign hamming[966] = 8'b11111111;
assign hamming[967] = 8'b10111001;
assign hamming[968] = 8'b00111000;
assign hamming[969] = 8'b00101000;
assign hamming[970] = 8'b00011000;
assign hamming[971] = 8'b01111000;
assign hamming[972] = 8'b01111001;
assign hamming[973] = 8'b00011001;
assign hamming[974] = 8'b00101001;
assign hamming[975] = 8'b00111001;
assign hamming[976] = 8'b00101010;
assign hamming[977] = 8'b00111010;
assign hamming[978] = 8'b01111010;
assign hamming[979] = 8'b00011010;
assign hamming[980] = 8'b00011011;
assign hamming[981] = 8'b01111011;
assign hamming[982] = 8'b00111011;
assign hamming[983] = 8'b00101011;
assign hamming[984] = 8'b11111111;
assign hamming[985] = 8'b10111010;
assign hamming[986] = 8'b11111111;
assign hamming[987] = 8'b11111111;
assign hamming[988] = 8'b11111111;
assign hamming[989] = 8'b11111111;
assign hamming[990] = 8'b10111011;
assign hamming[991] = 8'b11111111;
assign hamming[992] = 8'b00011100;
assign hamming[993] = 8'b01111100;
assign hamming[994] = 8'b00111100;
assign hamming[995] = 8'b00101100;
assign hamming[996] = 8'b00101101;
assign hamming[997] = 8'b00111101;
assign hamming[998] = 8'b01111101;
assign hamming[999] = 8'b00011101;
assign hamming[1000] = 8'b11111111;
assign hamming[1001] = 8'b11111111;
assign hamming[1002] = 8'b10111100;
assign hamming[1003] = 8'b11111111;
assign hamming[1004] = 8'b11111111;
assign hamming[1005] = 8'b10111101;
assign hamming[1006] = 8'b11111111;
assign hamming[1007] = 8'b11111111;
assign hamming[1008] = 8'b11111111;
assign hamming[1009] = 8'b11111111;
assign hamming[1010] = 8'b11111111;
assign hamming[1011] = 8'b10111110;
assign hamming[1012] = 8'b10111111;
assign hamming[1013] = 8'b11111111;
assign hamming[1014] = 8'b11111111;
assign hamming[1015] = 8'b11111111;
assign hamming[1016] = 8'b01111110;
assign hamming[1017] = 8'b00011110;
assign hamming[1018] = 8'b00101110;
assign hamming[1019] = 8'b00111110;
assign hamming[1020] = 8'b00111111;
assign hamming[1021] = 8'b00101111;
assign hamming[1022] = 8'b00011111;
assign hamming[1023] = 8'b01111111;
assign hamming[1024] = 8'b00000000;
assign hamming[1025] = 8'b01100000;
assign hamming[1026] = 8'b01010000;
assign hamming[1027] = 8'b01000000;
assign hamming[1028] = 8'b01000001;
assign hamming[1029] = 8'b01010001;
assign hamming[1030] = 8'b01100001;
assign hamming[1031] = 8'b00000001;
assign hamming[1032] = 8'b11111111;
assign hamming[1033] = 8'b11111111;
assign hamming[1034] = 8'b11111111;
assign hamming[1035] = 8'b11000000;
assign hamming[1036] = 8'b11000001;
assign hamming[1037] = 8'b11111111;
assign hamming[1038] = 8'b11111111;
assign hamming[1039] = 8'b11111111;
assign hamming[1040] = 8'b11111111;
assign hamming[1041] = 8'b11111111;
assign hamming[1042] = 8'b11000010;
assign hamming[1043] = 8'b11111111;
assign hamming[1044] = 8'b11111111;
assign hamming[1045] = 8'b11000011;
assign hamming[1046] = 8'b11111111;
assign hamming[1047] = 8'b11111111;
assign hamming[1048] = 8'b01100010;
assign hamming[1049] = 8'b00000010;
assign hamming[1050] = 8'b01000010;
assign hamming[1051] = 8'b01010010;
assign hamming[1052] = 8'b01010011;
assign hamming[1053] = 8'b01000011;
assign hamming[1054] = 8'b00000011;
assign hamming[1055] = 8'b01100011;
assign hamming[1056] = 8'b11111111;
assign hamming[1057] = 8'b11000100;
assign hamming[1058] = 8'b11111111;
assign hamming[1059] = 8'b11111111;
assign hamming[1060] = 8'b11111111;
assign hamming[1061] = 8'b11111111;
assign hamming[1062] = 8'b11000101;
assign hamming[1063] = 8'b11111111;
assign hamming[1064] = 8'b01010100;
assign hamming[1065] = 8'b01000100;
assign hamming[1066] = 8'b00000100;
assign hamming[1067] = 8'b01100100;
assign hamming[1068] = 8'b01100101;
assign hamming[1069] = 8'b00000101;
assign hamming[1070] = 8'b01000101;
assign hamming[1071] = 8'b01010101;
assign hamming[1072] = 8'b01000110;
assign hamming[1073] = 8'b01010110;
assign hamming[1074] = 8'b01100110;
assign hamming[1075] = 8'b00000110;
assign hamming[1076] = 8'b00000111;
assign hamming[1077] = 8'b01100111;
assign hamming[1078] = 8'b01010111;
assign hamming[1079] = 8'b01000111;
assign hamming[1080] = 8'b11000110;
assign hamming[1081] = 8'b11111111;
assign hamming[1082] = 8'b11111111;
assign hamming[1083] = 8'b11111111;
assign hamming[1084] = 8'b11111111;
assign hamming[1085] = 8'b11111111;
assign hamming[1086] = 8'b11111111;
assign hamming[1087] = 8'b11000111;
assign hamming[1088] = 8'b11001000;
assign hamming[1089] = 8'b11111111;
assign hamming[1090] = 8'b11111111;
assign hamming[1091] = 8'b11111111;
assign hamming[1092] = 8'b11111111;
assign hamming[1093] = 8'b11111111;
assign hamming[1094] = 8'b11111111;
assign hamming[1095] = 8'b11001001;
assign hamming[1096] = 8'b01001000;
assign hamming[1097] = 8'b01011000;
assign hamming[1098] = 8'b01101000;
assign hamming[1099] = 8'b00001000;
assign hamming[1100] = 8'b00001001;
assign hamming[1101] = 8'b01101001;
assign hamming[1102] = 8'b01011001;
assign hamming[1103] = 8'b01001001;
assign hamming[1104] = 8'b01011010;
assign hamming[1105] = 8'b01001010;
assign hamming[1106] = 8'b00001010;
assign hamming[1107] = 8'b01101010;
assign hamming[1108] = 8'b01101011;
assign hamming[1109] = 8'b00001011;
assign hamming[1110] = 8'b01001011;
assign hamming[1111] = 8'b01011011;
assign hamming[1112] = 8'b11111111;
assign hamming[1113] = 8'b11001010;
assign hamming[1114] = 8'b11111111;
assign hamming[1115] = 8'b11111111;
assign hamming[1116] = 8'b11111111;
assign hamming[1117] = 8'b11111111;
assign hamming[1118] = 8'b11001011;
assign hamming[1119] = 8'b11111111;
assign hamming[1120] = 8'b01101100;
assign hamming[1121] = 8'b00001100;
assign hamming[1122] = 8'b01001100;
assign hamming[1123] = 8'b01011100;
assign hamming[1124] = 8'b01011101;
assign hamming[1125] = 8'b01001101;
assign hamming[1126] = 8'b00001101;
assign hamming[1127] = 8'b01101101;
assign hamming[1128] = 8'b11111111;
assign hamming[1129] = 8'b11111111;
assign hamming[1130] = 8'b11001100;
assign hamming[1131] = 8'b11111111;
assign hamming[1132] = 8'b11111111;
assign hamming[1133] = 8'b11001101;
assign hamming[1134] = 8'b11111111;
assign hamming[1135] = 8'b11111111;
assign hamming[1136] = 8'b11111111;
assign hamming[1137] = 8'b11111111;
assign hamming[1138] = 8'b11111111;
assign hamming[1139] = 8'b11001110;
assign hamming[1140] = 8'b11001111;
assign hamming[1141] = 8'b11111111;
assign hamming[1142] = 8'b11111111;
assign hamming[1143] = 8'b11111111;
assign hamming[1144] = 8'b00001110;
assign hamming[1145] = 8'b01101110;
assign hamming[1146] = 8'b01011110;
assign hamming[1147] = 8'b01001110;
assign hamming[1148] = 8'b01001111;
assign hamming[1149] = 8'b01011111;
assign hamming[1150] = 8'b01101111;
assign hamming[1151] = 8'b00001111;
assign hamming[1152] = 8'b01000001;
assign hamming[1153] = 8'b01000000;
assign hamming[1154] = 8'b01000000;
assign hamming[1155] = 8'b01000000;
assign hamming[1156] = 8'b01000001;
assign hamming[1157] = 8'b01000001;
assign hamming[1158] = 8'b01000001;
assign hamming[1159] = 8'b01000000;
assign hamming[1160] = 8'b01001000;
assign hamming[1161] = 8'b01000100;
assign hamming[1162] = 8'b01000010;
assign hamming[1163] = 8'b01000000;
assign hamming[1164] = 8'b01000001;
assign hamming[1165] = 8'b01000011;
assign hamming[1166] = 8'b01000101;
assign hamming[1167] = 8'b01001001;
assign hamming[1168] = 8'b01000110;
assign hamming[1169] = 8'b01001010;
assign hamming[1170] = 8'b01000010;
assign hamming[1171] = 8'b01000000;
assign hamming[1172] = 8'b01000001;
assign hamming[1173] = 8'b01000011;
assign hamming[1174] = 8'b01001011;
assign hamming[1175] = 8'b01000111;
assign hamming[1176] = 8'b01000010;
assign hamming[1177] = 8'b01000011;
assign hamming[1178] = 8'b01000010;
assign hamming[1179] = 8'b01000010;
assign hamming[1180] = 8'b01000011;
assign hamming[1181] = 8'b01000011;
assign hamming[1182] = 8'b01000010;
assign hamming[1183] = 8'b01000011;
assign hamming[1184] = 8'b01000110;
assign hamming[1185] = 8'b01000100;
assign hamming[1186] = 8'b01001100;
assign hamming[1187] = 8'b01000000;
assign hamming[1188] = 8'b01000001;
assign hamming[1189] = 8'b01001101;
assign hamming[1190] = 8'b01000101;
assign hamming[1191] = 8'b01000111;
assign hamming[1192] = 8'b01000100;
assign hamming[1193] = 8'b01000100;
assign hamming[1194] = 8'b01000101;
assign hamming[1195] = 8'b01000100;
assign hamming[1196] = 8'b01000101;
assign hamming[1197] = 8'b01000100;
assign hamming[1198] = 8'b01000101;
assign hamming[1199] = 8'b01000101;
assign hamming[1200] = 8'b01000110;
assign hamming[1201] = 8'b01000110;
assign hamming[1202] = 8'b01000110;
assign hamming[1203] = 8'b01000111;
assign hamming[1204] = 8'b01000110;
assign hamming[1205] = 8'b01000111;
assign hamming[1206] = 8'b01000111;
assign hamming[1207] = 8'b01000111;
assign hamming[1208] = 8'b01000110;
assign hamming[1209] = 8'b01000100;
assign hamming[1210] = 8'b01000010;
assign hamming[1211] = 8'b01001110;
assign hamming[1212] = 8'b01001111;
assign hamming[1213] = 8'b01000011;
assign hamming[1214] = 8'b01000101;
assign hamming[1215] = 8'b01000111;
assign hamming[1216] = 8'b01001000;
assign hamming[1217] = 8'b01001010;
assign hamming[1218] = 8'b01001100;
assign hamming[1219] = 8'b01000000;
assign hamming[1220] = 8'b01000001;
assign hamming[1221] = 8'b01001101;
assign hamming[1222] = 8'b01001011;
assign hamming[1223] = 8'b01001001;
assign hamming[1224] = 8'b01001000;
assign hamming[1225] = 8'b01001000;
assign hamming[1226] = 8'b01001000;
assign hamming[1227] = 8'b01001001;
assign hamming[1228] = 8'b01001000;
assign hamming[1229] = 8'b01001001;
assign hamming[1230] = 8'b01001001;
assign hamming[1231] = 8'b01001001;
assign hamming[1232] = 8'b01001010;
assign hamming[1233] = 8'b01001010;
assign hamming[1234] = 8'b01001011;
assign hamming[1235] = 8'b01001010;
assign hamming[1236] = 8'b01001011;
assign hamming[1237] = 8'b01001010;
assign hamming[1238] = 8'b01001011;
assign hamming[1239] = 8'b01001011;
assign hamming[1240] = 8'b01001000;
assign hamming[1241] = 8'b01001010;
assign hamming[1242] = 8'b01000010;
assign hamming[1243] = 8'b01001110;
assign hamming[1244] = 8'b01001111;
assign hamming[1245] = 8'b01000011;
assign hamming[1246] = 8'b01001011;
assign hamming[1247] = 8'b01001001;
assign hamming[1248] = 8'b01001100;
assign hamming[1249] = 8'b01001101;
assign hamming[1250] = 8'b01001100;
assign hamming[1251] = 8'b01001100;
assign hamming[1252] = 8'b01001101;
assign hamming[1253] = 8'b01001101;
assign hamming[1254] = 8'b01001100;
assign hamming[1255] = 8'b01001101;
assign hamming[1256] = 8'b01001000;
assign hamming[1257] = 8'b01000100;
assign hamming[1258] = 8'b01001100;
assign hamming[1259] = 8'b01001110;
assign hamming[1260] = 8'b01001111;
assign hamming[1261] = 8'b01001101;
assign hamming[1262] = 8'b01000101;
assign hamming[1263] = 8'b01001001;
assign hamming[1264] = 8'b01000110;
assign hamming[1265] = 8'b01001010;
assign hamming[1266] = 8'b01001100;
assign hamming[1267] = 8'b01001110;
assign hamming[1268] = 8'b01001111;
assign hamming[1269] = 8'b01001101;
assign hamming[1270] = 8'b01001011;
assign hamming[1271] = 8'b01000111;
assign hamming[1272] = 8'b01001111;
assign hamming[1273] = 8'b01001110;
assign hamming[1274] = 8'b01001110;
assign hamming[1275] = 8'b01001110;
assign hamming[1276] = 8'b01001111;
assign hamming[1277] = 8'b01001111;
assign hamming[1278] = 8'b01001111;
assign hamming[1279] = 8'b01001110;
assign hamming[1280] = 8'b01010000;
assign hamming[1281] = 8'b01010001;
assign hamming[1282] = 8'b01010000;
assign hamming[1283] = 8'b01010000;
assign hamming[1284] = 8'b01010001;
assign hamming[1285] = 8'b01010001;
assign hamming[1286] = 8'b01010000;
assign hamming[1287] = 8'b01010001;
assign hamming[1288] = 8'b01010100;
assign hamming[1289] = 8'b01011000;
assign hamming[1290] = 8'b01010000;
assign hamming[1291] = 8'b01010010;
assign hamming[1292] = 8'b01010011;
assign hamming[1293] = 8'b01010001;
assign hamming[1294] = 8'b01011001;
assign hamming[1295] = 8'b01010101;
assign hamming[1296] = 8'b01011010;
assign hamming[1297] = 8'b01010110;
assign hamming[1298] = 8'b01010000;
assign hamming[1299] = 8'b01010010;
assign hamming[1300] = 8'b01010011;
assign hamming[1301] = 8'b01010001;
assign hamming[1302] = 8'b01010111;
assign hamming[1303] = 8'b01011011;
assign hamming[1304] = 8'b01010011;
assign hamming[1305] = 8'b01010010;
assign hamming[1306] = 8'b01010010;
assign hamming[1307] = 8'b01010010;
assign hamming[1308] = 8'b01010011;
assign hamming[1309] = 8'b01010011;
assign hamming[1310] = 8'b01010011;
assign hamming[1311] = 8'b01010010;
assign hamming[1312] = 8'b01010100;
assign hamming[1313] = 8'b01010110;
assign hamming[1314] = 8'b01010000;
assign hamming[1315] = 8'b01011100;
assign hamming[1316] = 8'b01011101;
assign hamming[1317] = 8'b01010001;
assign hamming[1318] = 8'b01010111;
assign hamming[1319] = 8'b01010101;
assign hamming[1320] = 8'b01010100;
assign hamming[1321] = 8'b01010100;
assign hamming[1322] = 8'b01010100;
assign hamming[1323] = 8'b01010101;
assign hamming[1324] = 8'b01010100;
assign hamming[1325] = 8'b01010101;
assign hamming[1326] = 8'b01010101;
assign hamming[1327] = 8'b01010101;
assign hamming[1328] = 8'b01010110;
assign hamming[1329] = 8'b01010110;
assign hamming[1330] = 8'b01010111;
assign hamming[1331] = 8'b01010110;
assign hamming[1332] = 8'b01010111;
assign hamming[1333] = 8'b01010110;
assign hamming[1334] = 8'b01010111;
assign hamming[1335] = 8'b01010111;
assign hamming[1336] = 8'b01010100;
assign hamming[1337] = 8'b01010110;
assign hamming[1338] = 8'b01011110;
assign hamming[1339] = 8'b01010010;
assign hamming[1340] = 8'b01010011;
assign hamming[1341] = 8'b01011111;
assign hamming[1342] = 8'b01010111;
assign hamming[1343] = 8'b01010101;
assign hamming[1344] = 8'b01011010;
assign hamming[1345] = 8'b01011000;
assign hamming[1346] = 8'b01010000;
assign hamming[1347] = 8'b01011100;
assign hamming[1348] = 8'b01011101;
assign hamming[1349] = 8'b01010001;
assign hamming[1350] = 8'b01011001;
assign hamming[1351] = 8'b01011011;
assign hamming[1352] = 8'b01011000;
assign hamming[1353] = 8'b01011000;
assign hamming[1354] = 8'b01011001;
assign hamming[1355] = 8'b01011000;
assign hamming[1356] = 8'b01011001;
assign hamming[1357] = 8'b01011000;
assign hamming[1358] = 8'b01011001;
assign hamming[1359] = 8'b01011001;
assign hamming[1360] = 8'b01011010;
assign hamming[1361] = 8'b01011010;
assign hamming[1362] = 8'b01011010;
assign hamming[1363] = 8'b01011011;
assign hamming[1364] = 8'b01011010;
assign hamming[1365] = 8'b01011011;
assign hamming[1366] = 8'b01011011;
assign hamming[1367] = 8'b01011011;
assign hamming[1368] = 8'b01011010;
assign hamming[1369] = 8'b01011000;
assign hamming[1370] = 8'b01011110;
assign hamming[1371] = 8'b01010010;
assign hamming[1372] = 8'b01010011;
assign hamming[1373] = 8'b01011111;
assign hamming[1374] = 8'b01011001;
assign hamming[1375] = 8'b01011011;
assign hamming[1376] = 8'b01011101;
assign hamming[1377] = 8'b01011100;
assign hamming[1378] = 8'b01011100;
assign hamming[1379] = 8'b01011100;
assign hamming[1380] = 8'b01011101;
assign hamming[1381] = 8'b01011101;
assign hamming[1382] = 8'b01011101;
assign hamming[1383] = 8'b01011100;
assign hamming[1384] = 8'b01010100;
assign hamming[1385] = 8'b01011000;
assign hamming[1386] = 8'b01011110;
assign hamming[1387] = 8'b01011100;
assign hamming[1388] = 8'b01011101;
assign hamming[1389] = 8'b01011111;
assign hamming[1390] = 8'b01011001;
assign hamming[1391] = 8'b01010101;
assign hamming[1392] = 8'b01011010;
assign hamming[1393] = 8'b01010110;
assign hamming[1394] = 8'b01011110;
assign hamming[1395] = 8'b01011100;
assign hamming[1396] = 8'b01011101;
assign hamming[1397] = 8'b01011111;
assign hamming[1398] = 8'b01010111;
assign hamming[1399] = 8'b01011011;
assign hamming[1400] = 8'b01011110;
assign hamming[1401] = 8'b01011111;
assign hamming[1402] = 8'b01011110;
assign hamming[1403] = 8'b01011110;
assign hamming[1404] = 8'b01011111;
assign hamming[1405] = 8'b01011111;
assign hamming[1406] = 8'b01011110;
assign hamming[1407] = 8'b01011111;
assign hamming[1408] = 8'b01110000;
assign hamming[1409] = 8'b00010000;
assign hamming[1410] = 8'b01010000;
assign hamming[1411] = 8'b01000000;
assign hamming[1412] = 8'b01000001;
assign hamming[1413] = 8'b01010001;
assign hamming[1414] = 8'b00010001;
assign hamming[1415] = 8'b01110001;
assign hamming[1416] = 8'b11111111;
assign hamming[1417] = 8'b11111111;
assign hamming[1418] = 8'b11010000;
assign hamming[1419] = 8'b11111111;
assign hamming[1420] = 8'b11111111;
assign hamming[1421] = 8'b11010001;
assign hamming[1422] = 8'b11111111;
assign hamming[1423] = 8'b11111111;
assign hamming[1424] = 8'b11111111;
assign hamming[1425] = 8'b11111111;
assign hamming[1426] = 8'b11111111;
assign hamming[1427] = 8'b11010010;
assign hamming[1428] = 8'b11010011;
assign hamming[1429] = 8'b11111111;
assign hamming[1430] = 8'b11111111;
assign hamming[1431] = 8'b11111111;
assign hamming[1432] = 8'b00010010;
assign hamming[1433] = 8'b01110010;
assign hamming[1434] = 8'b01000010;
assign hamming[1435] = 8'b01010010;
assign hamming[1436] = 8'b01010011;
assign hamming[1437] = 8'b01000011;
assign hamming[1438] = 8'b01110011;
assign hamming[1439] = 8'b00010011;
assign hamming[1440] = 8'b11010100;
assign hamming[1441] = 8'b11111111;
assign hamming[1442] = 8'b11111111;
assign hamming[1443] = 8'b11111111;
assign hamming[1444] = 8'b11111111;
assign hamming[1445] = 8'b11111111;
assign hamming[1446] = 8'b11111111;
assign hamming[1447] = 8'b11010101;
assign hamming[1448] = 8'b01010100;
assign hamming[1449] = 8'b01000100;
assign hamming[1450] = 8'b01110100;
assign hamming[1451] = 8'b00010100;
assign hamming[1452] = 8'b00010101;
assign hamming[1453] = 8'b01110101;
assign hamming[1454] = 8'b01000101;
assign hamming[1455] = 8'b01010101;
assign hamming[1456] = 8'b01000110;
assign hamming[1457] = 8'b01010110;
assign hamming[1458] = 8'b00010110;
assign hamming[1459] = 8'b01110110;
assign hamming[1460] = 8'b01110111;
assign hamming[1461] = 8'b00010111;
assign hamming[1462] = 8'b01010111;
assign hamming[1463] = 8'b01000111;
assign hamming[1464] = 8'b11111111;
assign hamming[1465] = 8'b11010110;
assign hamming[1466] = 8'b11111111;
assign hamming[1467] = 8'b11111111;
assign hamming[1468] = 8'b11111111;
assign hamming[1469] = 8'b11111111;
assign hamming[1470] = 8'b11010111;
assign hamming[1471] = 8'b11111111;
assign hamming[1472] = 8'b11111111;
assign hamming[1473] = 8'b11011000;
assign hamming[1474] = 8'b11111111;
assign hamming[1475] = 8'b11111111;
assign hamming[1476] = 8'b11111111;
assign hamming[1477] = 8'b11111111;
assign hamming[1478] = 8'b11011001;
assign hamming[1479] = 8'b11111111;
assign hamming[1480] = 8'b01001000;
assign hamming[1481] = 8'b01011000;
assign hamming[1482] = 8'b00011000;
assign hamming[1483] = 8'b01111000;
assign hamming[1484] = 8'b01111001;
assign hamming[1485] = 8'b00011001;
assign hamming[1486] = 8'b01011001;
assign hamming[1487] = 8'b01001001;
assign hamming[1488] = 8'b01011010;
assign hamming[1489] = 8'b01001010;
assign hamming[1490] = 8'b01111010;
assign hamming[1491] = 8'b00011010;
assign hamming[1492] = 8'b00011011;
assign hamming[1493] = 8'b01111011;
assign hamming[1494] = 8'b01001011;
assign hamming[1495] = 8'b01011011;
assign hamming[1496] = 8'b11011010;
assign hamming[1497] = 8'b11111111;
assign hamming[1498] = 8'b11111111;
assign hamming[1499] = 8'b11111111;
assign hamming[1500] = 8'b11111111;
assign hamming[1501] = 8'b11111111;
assign hamming[1502] = 8'b11111111;
assign hamming[1503] = 8'b11011011;
assign hamming[1504] = 8'b00011100;
assign hamming[1505] = 8'b01111100;
assign hamming[1506] = 8'b01001100;
assign hamming[1507] = 8'b01011100;
assign hamming[1508] = 8'b01011101;
assign hamming[1509] = 8'b01001101;
assign hamming[1510] = 8'b01111101;
assign hamming[1511] = 8'b00011101;
assign hamming[1512] = 8'b11111111;
assign hamming[1513] = 8'b11111111;
assign hamming[1514] = 8'b11111111;
assign hamming[1515] = 8'b11011100;
assign hamming[1516] = 8'b11011101;
assign hamming[1517] = 8'b11111111;
assign hamming[1518] = 8'b11111111;
assign hamming[1519] = 8'b11111111;
assign hamming[1520] = 8'b11111111;
assign hamming[1521] = 8'b11111111;
assign hamming[1522] = 8'b11011110;
assign hamming[1523] = 8'b11111111;
assign hamming[1524] = 8'b11111111;
assign hamming[1525] = 8'b11011111;
assign hamming[1526] = 8'b11111111;
assign hamming[1527] = 8'b11111111;
assign hamming[1528] = 8'b01111110;
assign hamming[1529] = 8'b00011110;
assign hamming[1530] = 8'b01011110;
assign hamming[1531] = 8'b01001110;
assign hamming[1532] = 8'b01001111;
assign hamming[1533] = 8'b01011111;
assign hamming[1534] = 8'b00011111;
assign hamming[1535] = 8'b01111111;
assign hamming[1536] = 8'b01100000;
assign hamming[1537] = 8'b01100000;
assign hamming[1538] = 8'b01100001;
assign hamming[1539] = 8'b01100000;
assign hamming[1540] = 8'b01100001;
assign hamming[1541] = 8'b01100000;
assign hamming[1542] = 8'b01100001;
assign hamming[1543] = 8'b01100001;
assign hamming[1544] = 8'b01100010;
assign hamming[1545] = 8'b01100000;
assign hamming[1546] = 8'b01101000;
assign hamming[1547] = 8'b01100100;
assign hamming[1548] = 8'b01100101;
assign hamming[1549] = 8'b01101001;
assign hamming[1550] = 8'b01100001;
assign hamming[1551] = 8'b01100011;
assign hamming[1552] = 8'b01100010;
assign hamming[1553] = 8'b01100000;
assign hamming[1554] = 8'b01100110;
assign hamming[1555] = 8'b01101010;
assign hamming[1556] = 8'b01101011;
assign hamming[1557] = 8'b01100111;
assign hamming[1558] = 8'b01100001;
assign hamming[1559] = 8'b01100011;
assign hamming[1560] = 8'b01100010;
assign hamming[1561] = 8'b01100010;
assign hamming[1562] = 8'b01100010;
assign hamming[1563] = 8'b01100011;
assign hamming[1564] = 8'b01100010;
assign hamming[1565] = 8'b01100011;
assign hamming[1566] = 8'b01100011;
assign hamming[1567] = 8'b01100011;
assign hamming[1568] = 8'b01101100;
assign hamming[1569] = 8'b01100000;
assign hamming[1570] = 8'b01100110;
assign hamming[1571] = 8'b01100100;
assign hamming[1572] = 8'b01100101;
assign hamming[1573] = 8'b01100111;
assign hamming[1574] = 8'b01100001;
assign hamming[1575] = 8'b01101101;
assign hamming[1576] = 8'b01100101;
assign hamming[1577] = 8'b01100100;
assign hamming[1578] = 8'b01100100;
assign hamming[1579] = 8'b01100100;
assign hamming[1580] = 8'b01100101;
assign hamming[1581] = 8'b01100101;
assign hamming[1582] = 8'b01100101;
assign hamming[1583] = 8'b01100100;
assign hamming[1584] = 8'b01100110;
assign hamming[1585] = 8'b01100111;
assign hamming[1586] = 8'b01100110;
assign hamming[1587] = 8'b01100110;
assign hamming[1588] = 8'b01100111;
assign hamming[1589] = 8'b01100111;
assign hamming[1590] = 8'b01100110;
assign hamming[1591] = 8'b01100111;
assign hamming[1592] = 8'b01100010;
assign hamming[1593] = 8'b01101110;
assign hamming[1594] = 8'b01100110;
assign hamming[1595] = 8'b01100100;
assign hamming[1596] = 8'b01100101;
assign hamming[1597] = 8'b01100111;
assign hamming[1598] = 8'b01101111;
assign hamming[1599] = 8'b01100011;
assign hamming[1600] = 8'b01101100;
assign hamming[1601] = 8'b01100000;
assign hamming[1602] = 8'b01101000;
assign hamming[1603] = 8'b01101010;
assign hamming[1604] = 8'b01101011;
assign hamming[1605] = 8'b01101001;
assign hamming[1606] = 8'b01100001;
assign hamming[1607] = 8'b01101101;
assign hamming[1608] = 8'b01101000;
assign hamming[1609] = 8'b01101001;
assign hamming[1610] = 8'b01101000;
assign hamming[1611] = 8'b01101000;
assign hamming[1612] = 8'b01101001;
assign hamming[1613] = 8'b01101001;
assign hamming[1614] = 8'b01101000;
assign hamming[1615] = 8'b01101001;
assign hamming[1616] = 8'b01101011;
assign hamming[1617] = 8'b01101010;
assign hamming[1618] = 8'b01101010;
assign hamming[1619] = 8'b01101010;
assign hamming[1620] = 8'b01101011;
assign hamming[1621] = 8'b01101011;
assign hamming[1622] = 8'b01101011;
assign hamming[1623] = 8'b01101010;
assign hamming[1624] = 8'b01100010;
assign hamming[1625] = 8'b01101110;
assign hamming[1626] = 8'b01101000;
assign hamming[1627] = 8'b01101010;
assign hamming[1628] = 8'b01101011;
assign hamming[1629] = 8'b01101001;
assign hamming[1630] = 8'b01101111;
assign hamming[1631] = 8'b01100011;
assign hamming[1632] = 8'b01101100;
assign hamming[1633] = 8'b01101100;
assign hamming[1634] = 8'b01101100;
assign hamming[1635] = 8'b01101101;
assign hamming[1636] = 8'b01101100;
assign hamming[1637] = 8'b01101101;
assign hamming[1638] = 8'b01101101;
assign hamming[1639] = 8'b01101101;
assign hamming[1640] = 8'b01101100;
assign hamming[1641] = 8'b01101110;
assign hamming[1642] = 8'b01101000;
assign hamming[1643] = 8'b01100100;
assign hamming[1644] = 8'b01100101;
assign hamming[1645] = 8'b01101001;
assign hamming[1646] = 8'b01101111;
assign hamming[1647] = 8'b01101101;
assign hamming[1648] = 8'b01101100;
assign hamming[1649] = 8'b01101110;
assign hamming[1650] = 8'b01100110;
assign hamming[1651] = 8'b01101010;
assign hamming[1652] = 8'b01101011;
assign hamming[1653] = 8'b01100111;
assign hamming[1654] = 8'b01101111;
assign hamming[1655] = 8'b01101101;
assign hamming[1656] = 8'b01101110;
assign hamming[1657] = 8'b01101110;
assign hamming[1658] = 8'b01101111;
assign hamming[1659] = 8'b01101110;
assign hamming[1660] = 8'b01101111;
assign hamming[1661] = 8'b01101110;
assign hamming[1662] = 8'b01101111;
assign hamming[1663] = 8'b01101111;
assign hamming[1664] = 8'b01110000;
assign hamming[1665] = 8'b01100000;
assign hamming[1666] = 8'b00100000;
assign hamming[1667] = 8'b01000000;
assign hamming[1668] = 8'b01000001;
assign hamming[1669] = 8'b00100001;
assign hamming[1670] = 8'b01100001;
assign hamming[1671] = 8'b01110001;
assign hamming[1672] = 8'b11111111;
assign hamming[1673] = 8'b11100000;
assign hamming[1674] = 8'b11111111;
assign hamming[1675] = 8'b11111111;
assign hamming[1676] = 8'b11111111;
assign hamming[1677] = 8'b11111111;
assign hamming[1678] = 8'b11100001;
assign hamming[1679] = 8'b11111111;
assign hamming[1680] = 8'b11100010;
assign hamming[1681] = 8'b11111111;
assign hamming[1682] = 8'b11111111;
assign hamming[1683] = 8'b11111111;
assign hamming[1684] = 8'b11111111;
assign hamming[1685] = 8'b11111111;
assign hamming[1686] = 8'b11111111;
assign hamming[1687] = 8'b11100011;
assign hamming[1688] = 8'b01100010;
assign hamming[1689] = 8'b01110010;
assign hamming[1690] = 8'b01000010;
assign hamming[1691] = 8'b00100010;
assign hamming[1692] = 8'b00100011;
assign hamming[1693] = 8'b01000011;
assign hamming[1694] = 8'b01110011;
assign hamming[1695] = 8'b01100011;
assign hamming[1696] = 8'b11111111;
assign hamming[1697] = 8'b11111111;
assign hamming[1698] = 8'b11111111;
assign hamming[1699] = 8'b11100100;
assign hamming[1700] = 8'b11100101;
assign hamming[1701] = 8'b11111111;
assign hamming[1702] = 8'b11111111;
assign hamming[1703] = 8'b11111111;
assign hamming[1704] = 8'b00100100;
assign hamming[1705] = 8'b01000100;
assign hamming[1706] = 8'b01110100;
assign hamming[1707] = 8'b01100100;
assign hamming[1708] = 8'b01100101;
assign hamming[1709] = 8'b01110101;
assign hamming[1710] = 8'b01000101;
assign hamming[1711] = 8'b00100101;
assign hamming[1712] = 8'b01000110;
assign hamming[1713] = 8'b00100110;
assign hamming[1714] = 8'b01100110;
assign hamming[1715] = 8'b01110110;
assign hamming[1716] = 8'b01110111;
assign hamming[1717] = 8'b01100111;
assign hamming[1718] = 8'b00100111;
assign hamming[1719] = 8'b01000111;
assign hamming[1720] = 8'b11111111;
assign hamming[1721] = 8'b11111111;
assign hamming[1722] = 8'b11100110;
assign hamming[1723] = 8'b11111111;
assign hamming[1724] = 8'b11111111;
assign hamming[1725] = 8'b11100111;
assign hamming[1726] = 8'b11111111;
assign hamming[1727] = 8'b11111111;
assign hamming[1728] = 8'b11111111;
assign hamming[1729] = 8'b11111111;
assign hamming[1730] = 8'b11101000;
assign hamming[1731] = 8'b11111111;
assign hamming[1732] = 8'b11111111;
assign hamming[1733] = 8'b11101001;
assign hamming[1734] = 8'b11111111;
assign hamming[1735] = 8'b11111111;
assign hamming[1736] = 8'b01001000;
assign hamming[1737] = 8'b00101000;
assign hamming[1738] = 8'b01101000;
assign hamming[1739] = 8'b01111000;
assign hamming[1740] = 8'b01111001;
assign hamming[1741] = 8'b01101001;
assign hamming[1742] = 8'b00101001;
assign hamming[1743] = 8'b01001001;
assign hamming[1744] = 8'b00101010;
assign hamming[1745] = 8'b01001010;
assign hamming[1746] = 8'b01111010;
assign hamming[1747] = 8'b01101010;
assign hamming[1748] = 8'b01101011;
assign hamming[1749] = 8'b01111011;
assign hamming[1750] = 8'b01001011;
assign hamming[1751] = 8'b00101011;
assign hamming[1752] = 8'b11111111;
assign hamming[1753] = 8'b11111111;
assign hamming[1754] = 8'b11111111;
assign hamming[1755] = 8'b11101010;
assign hamming[1756] = 8'b11101011;
assign hamming[1757] = 8'b11111111;
assign hamming[1758] = 8'b11111111;
assign hamming[1759] = 8'b11111111;
assign hamming[1760] = 8'b01101100;
assign hamming[1761] = 8'b01111100;
assign hamming[1762] = 8'b01001100;
assign hamming[1763] = 8'b00101100;
assign hamming[1764] = 8'b00101101;
assign hamming[1765] = 8'b01001101;
assign hamming[1766] = 8'b01111101;
assign hamming[1767] = 8'b01101101;
assign hamming[1768] = 8'b11101100;
assign hamming[1769] = 8'b11111111;
assign hamming[1770] = 8'b11111111;
assign hamming[1771] = 8'b11111111;
assign hamming[1772] = 8'b11111111;
assign hamming[1773] = 8'b11111111;
assign hamming[1774] = 8'b11111111;
assign hamming[1775] = 8'b11101101;
assign hamming[1776] = 8'b11111111;
assign hamming[1777] = 8'b11101110;
assign hamming[1778] = 8'b11111111;
assign hamming[1779] = 8'b11111111;
assign hamming[1780] = 8'b11111111;
assign hamming[1781] = 8'b11111111;
assign hamming[1782] = 8'b11101111;
assign hamming[1783] = 8'b11111111;
assign hamming[1784] = 8'b01111110;
assign hamming[1785] = 8'b01101110;
assign hamming[1786] = 8'b00101110;
assign hamming[1787] = 8'b01001110;
assign hamming[1788] = 8'b01001111;
assign hamming[1789] = 8'b00101111;
assign hamming[1790] = 8'b01101111;
assign hamming[1791] = 8'b01111111;
assign hamming[1792] = 8'b01110000;
assign hamming[1793] = 8'b01100000;
assign hamming[1794] = 8'b01010000;
assign hamming[1795] = 8'b00110000;
assign hamming[1796] = 8'b00110001;
assign hamming[1797] = 8'b01010001;
assign hamming[1798] = 8'b01100001;
assign hamming[1799] = 8'b01110001;
assign hamming[1800] = 8'b11110000;
assign hamming[1801] = 8'b11111111;
assign hamming[1802] = 8'b11111111;
assign hamming[1803] = 8'b11111111;
assign hamming[1804] = 8'b11111111;
assign hamming[1805] = 8'b11111111;
assign hamming[1806] = 8'b11111111;
assign hamming[1807] = 8'b11110001;
assign hamming[1808] = 8'b11111111;
assign hamming[1809] = 8'b11110010;
assign hamming[1810] = 8'b11111111;
assign hamming[1811] = 8'b11111111;
assign hamming[1812] = 8'b11111111;
assign hamming[1813] = 8'b11111111;
assign hamming[1814] = 8'b11110011;
assign hamming[1815] = 8'b11111111;
assign hamming[1816] = 8'b01100010;
assign hamming[1817] = 8'b01110010;
assign hamming[1818] = 8'b00110010;
assign hamming[1819] = 8'b01010010;
assign hamming[1820] = 8'b01010011;
assign hamming[1821] = 8'b00110011;
assign hamming[1822] = 8'b01110011;
assign hamming[1823] = 8'b01100011;
assign hamming[1824] = 8'b11111111;
assign hamming[1825] = 8'b11111111;
assign hamming[1826] = 8'b11110100;
assign hamming[1827] = 8'b11111111;
assign hamming[1828] = 8'b11111111;
assign hamming[1829] = 8'b11110101;
assign hamming[1830] = 8'b11111111;
assign hamming[1831] = 8'b11111111;
assign hamming[1832] = 8'b01010100;
assign hamming[1833] = 8'b00110100;
assign hamming[1834] = 8'b01110100;
assign hamming[1835] = 8'b01100100;
assign hamming[1836] = 8'b01100101;
assign hamming[1837] = 8'b01110101;
assign hamming[1838] = 8'b00110101;
assign hamming[1839] = 8'b01010101;
assign hamming[1840] = 8'b00110110;
assign hamming[1841] = 8'b01010110;
assign hamming[1842] = 8'b01100110;
assign hamming[1843] = 8'b01110110;
assign hamming[1844] = 8'b01110111;
assign hamming[1845] = 8'b01100111;
assign hamming[1846] = 8'b01010111;
assign hamming[1847] = 8'b00110111;
assign hamming[1848] = 8'b11111111;
assign hamming[1849] = 8'b11111111;
assign hamming[1850] = 8'b11111111;
assign hamming[1851] = 8'b11110110;
assign hamming[1852] = 8'b11110111;
assign hamming[1853] = 8'b11111111;
assign hamming[1854] = 8'b11111111;
assign hamming[1855] = 8'b11111111;
assign hamming[1856] = 8'b11111111;
assign hamming[1857] = 8'b11111111;
assign hamming[1858] = 8'b11111111;
assign hamming[1859] = 8'b11111000;
assign hamming[1860] = 8'b11111001;
assign hamming[1861] = 8'b11111111;
assign hamming[1862] = 8'b11111111;
assign hamming[1863] = 8'b11111111;
assign hamming[1864] = 8'b00111000;
assign hamming[1865] = 8'b01011000;
assign hamming[1866] = 8'b01101000;
assign hamming[1867] = 8'b01111000;
assign hamming[1868] = 8'b01111001;
assign hamming[1869] = 8'b01101001;
assign hamming[1870] = 8'b01011001;
assign hamming[1871] = 8'b00111001;
assign hamming[1872] = 8'b01011010;
assign hamming[1873] = 8'b00111010;
assign hamming[1874] = 8'b01111010;
assign hamming[1875] = 8'b01101010;
assign hamming[1876] = 8'b01101011;
assign hamming[1877] = 8'b01111011;
assign hamming[1878] = 8'b00111011;
assign hamming[1879] = 8'b01011011;
assign hamming[1880] = 8'b11111111;
assign hamming[1881] = 8'b11111111;
assign hamming[1882] = 8'b11111010;
assign hamming[1883] = 8'b11111111;
assign hamming[1884] = 8'b11111111;
assign hamming[1885] = 8'b11111011;
assign hamming[1886] = 8'b11111111;
assign hamming[1887] = 8'b11111111;
assign hamming[1888] = 8'b01101100;
assign hamming[1889] = 8'b01111100;
assign hamming[1890] = 8'b00111100;
assign hamming[1891] = 8'b01011100;
assign hamming[1892] = 8'b01011101;
assign hamming[1893] = 8'b00111101;
assign hamming[1894] = 8'b01111101;
assign hamming[1895] = 8'b01101101;
assign hamming[1896] = 8'b11111111;
assign hamming[1897] = 8'b11111100;
assign hamming[1898] = 8'b11111111;
assign hamming[1899] = 8'b11111111;
assign hamming[1900] = 8'b11111111;
assign hamming[1901] = 8'b11111111;
assign hamming[1902] = 8'b11111101;
assign hamming[1903] = 8'b11111111;
assign hamming[1904] = 8'b11111110;
assign hamming[1905] = 8'b11111111;
assign hamming[1906] = 8'b11111111;
assign hamming[1907] = 8'b11111111;
assign hamming[1908] = 8'b11111111;
assign hamming[1909] = 8'b11111111;
assign hamming[1910] = 8'b11111111;
assign hamming[1911] = 8'b11111111;
assign hamming[1912] = 8'b01111110;
assign hamming[1913] = 8'b01101110;
assign hamming[1914] = 8'b01011110;
assign hamming[1915] = 8'b00111110;
assign hamming[1916] = 8'b00111111;
assign hamming[1917] = 8'b01011111;
assign hamming[1918] = 8'b01101111;
assign hamming[1919] = 8'b01111111;
assign hamming[1920] = 8'b01110000;
assign hamming[1921] = 8'b01110000;
assign hamming[1922] = 8'b01110000;
assign hamming[1923] = 8'b01110001;
assign hamming[1924] = 8'b01110000;
assign hamming[1925] = 8'b01110001;
assign hamming[1926] = 8'b01110001;
assign hamming[1927] = 8'b01110001;
assign hamming[1928] = 8'b01110000;
assign hamming[1929] = 8'b01110010;
assign hamming[1930] = 8'b01110100;
assign hamming[1931] = 8'b01111000;
assign hamming[1932] = 8'b01111001;
assign hamming[1933] = 8'b01110101;
assign hamming[1934] = 8'b01110011;
assign hamming[1935] = 8'b01110001;
assign hamming[1936] = 8'b01110000;
assign hamming[1937] = 8'b01110010;
assign hamming[1938] = 8'b01111010;
assign hamming[1939] = 8'b01110110;
assign hamming[1940] = 8'b01110111;
assign hamming[1941] = 8'b01111011;
assign hamming[1942] = 8'b01110011;
assign hamming[1943] = 8'b01110001;
assign hamming[1944] = 8'b01110010;
assign hamming[1945] = 8'b01110010;
assign hamming[1946] = 8'b01110011;
assign hamming[1947] = 8'b01110010;
assign hamming[1948] = 8'b01110011;
assign hamming[1949] = 8'b01110010;
assign hamming[1950] = 8'b01110011;
assign hamming[1951] = 8'b01110011;
assign hamming[1952] = 8'b01110000;
assign hamming[1953] = 8'b01111100;
assign hamming[1954] = 8'b01110100;
assign hamming[1955] = 8'b01110110;
assign hamming[1956] = 8'b01110111;
assign hamming[1957] = 8'b01110101;
assign hamming[1958] = 8'b01111101;
assign hamming[1959] = 8'b01110001;
assign hamming[1960] = 8'b01110100;
assign hamming[1961] = 8'b01110101;
assign hamming[1962] = 8'b01110100;
assign hamming[1963] = 8'b01110100;
assign hamming[1964] = 8'b01110101;
assign hamming[1965] = 8'b01110101;
assign hamming[1966] = 8'b01110100;
assign hamming[1967] = 8'b01110101;
assign hamming[1968] = 8'b01110111;
assign hamming[1969] = 8'b01110110;
assign hamming[1970] = 8'b01110110;
assign hamming[1971] = 8'b01110110;
assign hamming[1972] = 8'b01110111;
assign hamming[1973] = 8'b01110111;
assign hamming[1974] = 8'b01110111;
assign hamming[1975] = 8'b01110110;
assign hamming[1976] = 8'b01111110;
assign hamming[1977] = 8'b01110010;
assign hamming[1978] = 8'b01110100;
assign hamming[1979] = 8'b01110110;
assign hamming[1980] = 8'b01110111;
assign hamming[1981] = 8'b01110101;
assign hamming[1982] = 8'b01110011;
assign hamming[1983] = 8'b01111111;
assign hamming[1984] = 8'b01110000;
assign hamming[1985] = 8'b01111100;
assign hamming[1986] = 8'b01111010;
assign hamming[1987] = 8'b01111000;
assign hamming[1988] = 8'b01111001;
assign hamming[1989] = 8'b01111011;
assign hamming[1990] = 8'b01111101;
assign hamming[1991] = 8'b01110001;
assign hamming[1992] = 8'b01111001;
assign hamming[1993] = 8'b01111000;
assign hamming[1994] = 8'b01111000;
assign hamming[1995] = 8'b01111000;
assign hamming[1996] = 8'b01111001;
assign hamming[1997] = 8'b01111001;
assign hamming[1998] = 8'b01111001;
assign hamming[1999] = 8'b01111000;
assign hamming[2000] = 8'b01111010;
assign hamming[2001] = 8'b01111011;
assign hamming[2002] = 8'b01111010;
assign hamming[2003] = 8'b01111010;
assign hamming[2004] = 8'b01111011;
assign hamming[2005] = 8'b01111011;
assign hamming[2006] = 8'b01111010;
assign hamming[2007] = 8'b01111011;
assign hamming[2008] = 8'b01111110;
assign hamming[2009] = 8'b01110010;
assign hamming[2010] = 8'b01111010;
assign hamming[2011] = 8'b01111000;
assign hamming[2012] = 8'b01111001;
assign hamming[2013] = 8'b01111011;
assign hamming[2014] = 8'b01110011;
assign hamming[2015] = 8'b01111111;
assign hamming[2016] = 8'b01111100;
assign hamming[2017] = 8'b01111100;
assign hamming[2018] = 8'b01111101;
assign hamming[2019] = 8'b01111100;
assign hamming[2020] = 8'b01111101;
assign hamming[2021] = 8'b01111100;
assign hamming[2022] = 8'b01111101;
assign hamming[2023] = 8'b01111101;
assign hamming[2024] = 8'b01111110;
assign hamming[2025] = 8'b01111100;
assign hamming[2026] = 8'b01110100;
assign hamming[2027] = 8'b01111000;
assign hamming[2028] = 8'b01111001;
assign hamming[2029] = 8'b01110101;
assign hamming[2030] = 8'b01111101;
assign hamming[2031] = 8'b01111111;
assign hamming[2032] = 8'b01111110;
assign hamming[2033] = 8'b01111100;
assign hamming[2034] = 8'b01111010;
assign hamming[2035] = 8'b01110110;
assign hamming[2036] = 8'b01110111;
assign hamming[2037] = 8'b01111011;
assign hamming[2038] = 8'b01111101;
assign hamming[2039] = 8'b01111111;
assign hamming[2040] = 8'b01111110;
assign hamming[2041] = 8'b01111110;
assign hamming[2042] = 8'b01111110;
assign hamming[2043] = 8'b01111111;
assign hamming[2044] = 8'b01111110;
assign hamming[2045] = 8'b01111111;
assign hamming[2046] = 8'b01111111;
assign hamming[2047] = 8'b01111111;
assign hamming[2048] = 8'b00000000;
assign hamming[2049] = 8'b11111111;
assign hamming[2050] = 8'b11111111;
assign hamming[2051] = 8'b11111111;
assign hamming[2052] = 8'b11111111;
assign hamming[2053] = 8'b11111111;
assign hamming[2054] = 8'b11111111;
assign hamming[2055] = 8'b00000001;
assign hamming[2056] = 8'b10000000;
assign hamming[2057] = 8'b10010000;
assign hamming[2058] = 8'b10100000;
assign hamming[2059] = 8'b11000000;
assign hamming[2060] = 8'b11000001;
assign hamming[2061] = 8'b10100001;
assign hamming[2062] = 8'b10010001;
assign hamming[2063] = 8'b10000001;
assign hamming[2064] = 8'b10010010;
assign hamming[2065] = 8'b10000010;
assign hamming[2066] = 8'b11000010;
assign hamming[2067] = 8'b10100010;
assign hamming[2068] = 8'b10100011;
assign hamming[2069] = 8'b11000011;
assign hamming[2070] = 8'b10000011;
assign hamming[2071] = 8'b10010011;
assign hamming[2072] = 8'b11111111;
assign hamming[2073] = 8'b00000010;
assign hamming[2074] = 8'b11111111;
assign hamming[2075] = 8'b11111111;
assign hamming[2076] = 8'b11111111;
assign hamming[2077] = 8'b11111111;
assign hamming[2078] = 8'b00000011;
assign hamming[2079] = 8'b11111111;
assign hamming[2080] = 8'b10100100;
assign hamming[2081] = 8'b11000100;
assign hamming[2082] = 8'b10000100;
assign hamming[2083] = 8'b10010100;
assign hamming[2084] = 8'b10010101;
assign hamming[2085] = 8'b10000101;
assign hamming[2086] = 8'b11000101;
assign hamming[2087] = 8'b10100101;
assign hamming[2088] = 8'b11111111;
assign hamming[2089] = 8'b11111111;
assign hamming[2090] = 8'b00000100;
assign hamming[2091] = 8'b11111111;
assign hamming[2092] = 8'b11111111;
assign hamming[2093] = 8'b00000101;
assign hamming[2094] = 8'b11111111;
assign hamming[2095] = 8'b11111111;
assign hamming[2096] = 8'b11111111;
assign hamming[2097] = 8'b11111111;
assign hamming[2098] = 8'b11111111;
assign hamming[2099] = 8'b00000110;
assign hamming[2100] = 8'b00000111;
assign hamming[2101] = 8'b11111111;
assign hamming[2102] = 8'b11111111;
assign hamming[2103] = 8'b11111111;
assign hamming[2104] = 8'b11000110;
assign hamming[2105] = 8'b10100110;
assign hamming[2106] = 8'b10010110;
assign hamming[2107] = 8'b10000110;
assign hamming[2108] = 8'b10000111;
assign hamming[2109] = 8'b10010111;
assign hamming[2110] = 8'b10100111;
assign hamming[2111] = 8'b11000111;
assign hamming[2112] = 8'b11001000;
assign hamming[2113] = 8'b10101000;
assign hamming[2114] = 8'b10011000;
assign hamming[2115] = 8'b10001000;
assign hamming[2116] = 8'b10001001;
assign hamming[2117] = 8'b10011001;
assign hamming[2118] = 8'b10101001;
assign hamming[2119] = 8'b11001001;
assign hamming[2120] = 8'b11111111;
assign hamming[2121] = 8'b11111111;
assign hamming[2122] = 8'b11111111;
assign hamming[2123] = 8'b00001000;
assign hamming[2124] = 8'b00001001;
assign hamming[2125] = 8'b11111111;
assign hamming[2126] = 8'b11111111;
assign hamming[2127] = 8'b11111111;
assign hamming[2128] = 8'b11111111;
assign hamming[2129] = 8'b11111111;
assign hamming[2130] = 8'b00001010;
assign hamming[2131] = 8'b11111111;
assign hamming[2132] = 8'b11111111;
assign hamming[2133] = 8'b00001011;
assign hamming[2134] = 8'b11111111;
assign hamming[2135] = 8'b11111111;
assign hamming[2136] = 8'b10101010;
assign hamming[2137] = 8'b11001010;
assign hamming[2138] = 8'b10001010;
assign hamming[2139] = 8'b10011010;
assign hamming[2140] = 8'b10011011;
assign hamming[2141] = 8'b10001011;
assign hamming[2142] = 8'b11001011;
assign hamming[2143] = 8'b10101011;
assign hamming[2144] = 8'b11111111;
assign hamming[2145] = 8'b00001100;
assign hamming[2146] = 8'b11111111;
assign hamming[2147] = 8'b11111111;
assign hamming[2148] = 8'b11111111;
assign hamming[2149] = 8'b11111111;
assign hamming[2150] = 8'b00001101;
assign hamming[2151] = 8'b11111111;
assign hamming[2152] = 8'b10011100;
assign hamming[2153] = 8'b10001100;
assign hamming[2154] = 8'b11001100;
assign hamming[2155] = 8'b10101100;
assign hamming[2156] = 8'b10101101;
assign hamming[2157] = 8'b11001101;
assign hamming[2158] = 8'b10001101;
assign hamming[2159] = 8'b10011101;
assign hamming[2160] = 8'b10001110;
assign hamming[2161] = 8'b10011110;
assign hamming[2162] = 8'b10101110;
assign hamming[2163] = 8'b11001110;
assign hamming[2164] = 8'b11001111;
assign hamming[2165] = 8'b10101111;
assign hamming[2166] = 8'b10011111;
assign hamming[2167] = 8'b10001111;
assign hamming[2168] = 8'b00001110;
assign hamming[2169] = 8'b11111111;
assign hamming[2170] = 8'b11111111;
assign hamming[2171] = 8'b11111111;
assign hamming[2172] = 8'b11111111;
assign hamming[2173] = 8'b11111111;
assign hamming[2174] = 8'b11111111;
assign hamming[2175] = 8'b00001111;
assign hamming[2176] = 8'b10000000;
assign hamming[2177] = 8'b10000010;
assign hamming[2178] = 8'b10000100;
assign hamming[2179] = 8'b10001000;
assign hamming[2180] = 8'b10001001;
assign hamming[2181] = 8'b10000101;
assign hamming[2182] = 8'b10000011;
assign hamming[2183] = 8'b10000001;
assign hamming[2184] = 8'b10000000;
assign hamming[2185] = 8'b10000000;
assign hamming[2186] = 8'b10000000;
assign hamming[2187] = 8'b10000001;
assign hamming[2188] = 8'b10000000;
assign hamming[2189] = 8'b10000001;
assign hamming[2190] = 8'b10000001;
assign hamming[2191] = 8'b10000001;
assign hamming[2192] = 8'b10000010;
assign hamming[2193] = 8'b10000010;
assign hamming[2194] = 8'b10000011;
assign hamming[2195] = 8'b10000010;
assign hamming[2196] = 8'b10000011;
assign hamming[2197] = 8'b10000010;
assign hamming[2198] = 8'b10000011;
assign hamming[2199] = 8'b10000011;
assign hamming[2200] = 8'b10000000;
assign hamming[2201] = 8'b10000010;
assign hamming[2202] = 8'b10001010;
assign hamming[2203] = 8'b10000110;
assign hamming[2204] = 8'b10000111;
assign hamming[2205] = 8'b10001011;
assign hamming[2206] = 8'b10000011;
assign hamming[2207] = 8'b10000001;
assign hamming[2208] = 8'b10000100;
assign hamming[2209] = 8'b10000101;
assign hamming[2210] = 8'b10000100;
assign hamming[2211] = 8'b10000100;
assign hamming[2212] = 8'b10000101;
assign hamming[2213] = 8'b10000101;
assign hamming[2214] = 8'b10000100;
assign hamming[2215] = 8'b10000101;
assign hamming[2216] = 8'b10000000;
assign hamming[2217] = 8'b10001100;
assign hamming[2218] = 8'b10000100;
assign hamming[2219] = 8'b10000110;
assign hamming[2220] = 8'b10000111;
assign hamming[2221] = 8'b10000101;
assign hamming[2222] = 8'b10001101;
assign hamming[2223] = 8'b10000001;
assign hamming[2224] = 8'b10001110;
assign hamming[2225] = 8'b10000010;
assign hamming[2226] = 8'b10000100;
assign hamming[2227] = 8'b10000110;
assign hamming[2228] = 8'b10000111;
assign hamming[2229] = 8'b10000101;
assign hamming[2230] = 8'b10000011;
assign hamming[2231] = 8'b10001111;
assign hamming[2232] = 8'b10000111;
assign hamming[2233] = 8'b10000110;
assign hamming[2234] = 8'b10000110;
assign hamming[2235] = 8'b10000110;
assign hamming[2236] = 8'b10000111;
assign hamming[2237] = 8'b10000111;
assign hamming[2238] = 8'b10000111;
assign hamming[2239] = 8'b10000110;
assign hamming[2240] = 8'b10001001;
assign hamming[2241] = 8'b10001000;
assign hamming[2242] = 8'b10001000;
assign hamming[2243] = 8'b10001000;
assign hamming[2244] = 8'b10001001;
assign hamming[2245] = 8'b10001001;
assign hamming[2246] = 8'b10001001;
assign hamming[2247] = 8'b10001000;
assign hamming[2248] = 8'b10000000;
assign hamming[2249] = 8'b10001100;
assign hamming[2250] = 8'b10001010;
assign hamming[2251] = 8'b10001000;
assign hamming[2252] = 8'b10001001;
assign hamming[2253] = 8'b10001011;
assign hamming[2254] = 8'b10001101;
assign hamming[2255] = 8'b10000001;
assign hamming[2256] = 8'b10001110;
assign hamming[2257] = 8'b10000010;
assign hamming[2258] = 8'b10001010;
assign hamming[2259] = 8'b10001000;
assign hamming[2260] = 8'b10001001;
assign hamming[2261] = 8'b10001011;
assign hamming[2262] = 8'b10000011;
assign hamming[2263] = 8'b10001111;
assign hamming[2264] = 8'b10001010;
assign hamming[2265] = 8'b10001011;
assign hamming[2266] = 8'b10001010;
assign hamming[2267] = 8'b10001010;
assign hamming[2268] = 8'b10001011;
assign hamming[2269] = 8'b10001011;
assign hamming[2270] = 8'b10001010;
assign hamming[2271] = 8'b10001011;
assign hamming[2272] = 8'b10001110;
assign hamming[2273] = 8'b10001100;
assign hamming[2274] = 8'b10000100;
assign hamming[2275] = 8'b10001000;
assign hamming[2276] = 8'b10001001;
assign hamming[2277] = 8'b10000101;
assign hamming[2278] = 8'b10001101;
assign hamming[2279] = 8'b10001111;
assign hamming[2280] = 8'b10001100;
assign hamming[2281] = 8'b10001100;
assign hamming[2282] = 8'b10001101;
assign hamming[2283] = 8'b10001100;
assign hamming[2284] = 8'b10001101;
assign hamming[2285] = 8'b10001100;
assign hamming[2286] = 8'b10001101;
assign hamming[2287] = 8'b10001101;
assign hamming[2288] = 8'b10001110;
assign hamming[2289] = 8'b10001110;
assign hamming[2290] = 8'b10001110;
assign hamming[2291] = 8'b10001111;
assign hamming[2292] = 8'b10001110;
assign hamming[2293] = 8'b10001111;
assign hamming[2294] = 8'b10001111;
assign hamming[2295] = 8'b10001111;
assign hamming[2296] = 8'b10001110;
assign hamming[2297] = 8'b10001100;
assign hamming[2298] = 8'b10001010;
assign hamming[2299] = 8'b10000110;
assign hamming[2300] = 8'b10000111;
assign hamming[2301] = 8'b10001011;
assign hamming[2302] = 8'b10001101;
assign hamming[2303] = 8'b10001111;
assign hamming[2304] = 8'b10010010;
assign hamming[2305] = 8'b10010000;
assign hamming[2306] = 8'b10011000;
assign hamming[2307] = 8'b10010100;
assign hamming[2308] = 8'b10010101;
assign hamming[2309] = 8'b10011001;
assign hamming[2310] = 8'b10010001;
assign hamming[2311] = 8'b10010011;
assign hamming[2312] = 8'b10010000;
assign hamming[2313] = 8'b10010000;
assign hamming[2314] = 8'b10010001;
assign hamming[2315] = 8'b10010000;
assign hamming[2316] = 8'b10010001;
assign hamming[2317] = 8'b10010000;
assign hamming[2318] = 8'b10010001;
assign hamming[2319] = 8'b10010001;
assign hamming[2320] = 8'b10010010;
assign hamming[2321] = 8'b10010010;
assign hamming[2322] = 8'b10010010;
assign hamming[2323] = 8'b10010011;
assign hamming[2324] = 8'b10010010;
assign hamming[2325] = 8'b10010011;
assign hamming[2326] = 8'b10010011;
assign hamming[2327] = 8'b10010011;
assign hamming[2328] = 8'b10010010;
assign hamming[2329] = 8'b10010000;
assign hamming[2330] = 8'b10010110;
assign hamming[2331] = 8'b10011010;
assign hamming[2332] = 8'b10011011;
assign hamming[2333] = 8'b10010111;
assign hamming[2334] = 8'b10010001;
assign hamming[2335] = 8'b10010011;
assign hamming[2336] = 8'b10010101;
assign hamming[2337] = 8'b10010100;
assign hamming[2338] = 8'b10010100;
assign hamming[2339] = 8'b10010100;
assign hamming[2340] = 8'b10010101;
assign hamming[2341] = 8'b10010101;
assign hamming[2342] = 8'b10010101;
assign hamming[2343] = 8'b10010100;
assign hamming[2344] = 8'b10011100;
assign hamming[2345] = 8'b10010000;
assign hamming[2346] = 8'b10010110;
assign hamming[2347] = 8'b10010100;
assign hamming[2348] = 8'b10010101;
assign hamming[2349] = 8'b10010111;
assign hamming[2350] = 8'b10010001;
assign hamming[2351] = 8'b10011101;
assign hamming[2352] = 8'b10010010;
assign hamming[2353] = 8'b10011110;
assign hamming[2354] = 8'b10010110;
assign hamming[2355] = 8'b10010100;
assign hamming[2356] = 8'b10010101;
assign hamming[2357] = 8'b10010111;
assign hamming[2358] = 8'b10011111;
assign hamming[2359] = 8'b10010011;
assign hamming[2360] = 8'b10010110;
assign hamming[2361] = 8'b10010111;
assign hamming[2362] = 8'b10010110;
assign hamming[2363] = 8'b10010110;
assign hamming[2364] = 8'b10010111;
assign hamming[2365] = 8'b10010111;
assign hamming[2366] = 8'b10010110;
assign hamming[2367] = 8'b10010111;
assign hamming[2368] = 8'b10011000;
assign hamming[2369] = 8'b10011001;
assign hamming[2370] = 8'b10011000;
assign hamming[2371] = 8'b10011000;
assign hamming[2372] = 8'b10011001;
assign hamming[2373] = 8'b10011001;
assign hamming[2374] = 8'b10011000;
assign hamming[2375] = 8'b10011001;
assign hamming[2376] = 8'b10011100;
assign hamming[2377] = 8'b10010000;
assign hamming[2378] = 8'b10011000;
assign hamming[2379] = 8'b10011010;
assign hamming[2380] = 8'b10011011;
assign hamming[2381] = 8'b10011001;
assign hamming[2382] = 8'b10010001;
assign hamming[2383] = 8'b10011101;
assign hamming[2384] = 8'b10010010;
assign hamming[2385] = 8'b10011110;
assign hamming[2386] = 8'b10011000;
assign hamming[2387] = 8'b10011010;
assign hamming[2388] = 8'b10011011;
assign hamming[2389] = 8'b10011001;
assign hamming[2390] = 8'b10011111;
assign hamming[2391] = 8'b10010011;
assign hamming[2392] = 8'b10011011;
assign hamming[2393] = 8'b10011010;
assign hamming[2394] = 8'b10011010;
assign hamming[2395] = 8'b10011010;
assign hamming[2396] = 8'b10011011;
assign hamming[2397] = 8'b10011011;
assign hamming[2398] = 8'b10011011;
assign hamming[2399] = 8'b10011010;
assign hamming[2400] = 8'b10011100;
assign hamming[2401] = 8'b10011110;
assign hamming[2402] = 8'b10011000;
assign hamming[2403] = 8'b10010100;
assign hamming[2404] = 8'b10010101;
assign hamming[2405] = 8'b10011001;
assign hamming[2406] = 8'b10011111;
assign hamming[2407] = 8'b10011101;
assign hamming[2408] = 8'b10011100;
assign hamming[2409] = 8'b10011100;
assign hamming[2410] = 8'b10011100;
assign hamming[2411] = 8'b10011101;
assign hamming[2412] = 8'b10011100;
assign hamming[2413] = 8'b10011101;
assign hamming[2414] = 8'b10011101;
assign hamming[2415] = 8'b10011101;
assign hamming[2416] = 8'b10011110;
assign hamming[2417] = 8'b10011110;
assign hamming[2418] = 8'b10011111;
assign hamming[2419] = 8'b10011110;
assign hamming[2420] = 8'b10011111;
assign hamming[2421] = 8'b10011110;
assign hamming[2422] = 8'b10011111;
assign hamming[2423] = 8'b10011111;
assign hamming[2424] = 8'b10011100;
assign hamming[2425] = 8'b10011110;
assign hamming[2426] = 8'b10010110;
assign hamming[2427] = 8'b10011010;
assign hamming[2428] = 8'b10011011;
assign hamming[2429] = 8'b10010111;
assign hamming[2430] = 8'b10011111;
assign hamming[2431] = 8'b10011101;
assign hamming[2432] = 8'b11111111;
assign hamming[2433] = 8'b00010000;
assign hamming[2434] = 8'b11111111;
assign hamming[2435] = 8'b11111111;
assign hamming[2436] = 8'b11111111;
assign hamming[2437] = 8'b11111111;
assign hamming[2438] = 8'b00010001;
assign hamming[2439] = 8'b11111111;
assign hamming[2440] = 8'b10000000;
assign hamming[2441] = 8'b10010000;
assign hamming[2442] = 8'b11010000;
assign hamming[2443] = 8'b10110000;
assign hamming[2444] = 8'b10110001;
assign hamming[2445] = 8'b11010001;
assign hamming[2446] = 8'b10010001;
assign hamming[2447] = 8'b10000001;
assign hamming[2448] = 8'b10010010;
assign hamming[2449] = 8'b10000010;
assign hamming[2450] = 8'b10110010;
assign hamming[2451] = 8'b11010010;
assign hamming[2452] = 8'b11010011;
assign hamming[2453] = 8'b10110011;
assign hamming[2454] = 8'b10000011;
assign hamming[2455] = 8'b10010011;
assign hamming[2456] = 8'b00010010;
assign hamming[2457] = 8'b11111111;
assign hamming[2458] = 8'b11111111;
assign hamming[2459] = 8'b11111111;
assign hamming[2460] = 8'b11111111;
assign hamming[2461] = 8'b11111111;
assign hamming[2462] = 8'b11111111;
assign hamming[2463] = 8'b00010011;
assign hamming[2464] = 8'b11010100;
assign hamming[2465] = 8'b10110100;
assign hamming[2466] = 8'b10000100;
assign hamming[2467] = 8'b10010100;
assign hamming[2468] = 8'b10010101;
assign hamming[2469] = 8'b10000101;
assign hamming[2470] = 8'b10110101;
assign hamming[2471] = 8'b11010101;
assign hamming[2472] = 8'b11111111;
assign hamming[2473] = 8'b11111111;
assign hamming[2474] = 8'b11111111;
assign hamming[2475] = 8'b00010100;
assign hamming[2476] = 8'b00010101;
assign hamming[2477] = 8'b11111111;
assign hamming[2478] = 8'b11111111;
assign hamming[2479] = 8'b11111111;
assign hamming[2480] = 8'b11111111;
assign hamming[2481] = 8'b11111111;
assign hamming[2482] = 8'b00010110;
assign hamming[2483] = 8'b11111111;
assign hamming[2484] = 8'b11111111;
assign hamming[2485] = 8'b00010111;
assign hamming[2486] = 8'b11111111;
assign hamming[2487] = 8'b11111111;
assign hamming[2488] = 8'b10110110;
assign hamming[2489] = 8'b11010110;
assign hamming[2490] = 8'b10010110;
assign hamming[2491] = 8'b10000110;
assign hamming[2492] = 8'b10000111;
assign hamming[2493] = 8'b10010111;
assign hamming[2494] = 8'b11010111;
assign hamming[2495] = 8'b10110111;
assign hamming[2496] = 8'b10111000;
assign hamming[2497] = 8'b11011000;
assign hamming[2498] = 8'b10011000;
assign hamming[2499] = 8'b10001000;
assign hamming[2500] = 8'b10001001;
assign hamming[2501] = 8'b10011001;
assign hamming[2502] = 8'b11011001;
assign hamming[2503] = 8'b10111001;
assign hamming[2504] = 8'b11111111;
assign hamming[2505] = 8'b11111111;
assign hamming[2506] = 8'b00011000;
assign hamming[2507] = 8'b11111111;
assign hamming[2508] = 8'b11111111;
assign hamming[2509] = 8'b00011001;
assign hamming[2510] = 8'b11111111;
assign hamming[2511] = 8'b11111111;
assign hamming[2512] = 8'b11111111;
assign hamming[2513] = 8'b11111111;
assign hamming[2514] = 8'b11111111;
assign hamming[2515] = 8'b00011010;
assign hamming[2516] = 8'b00011011;
assign hamming[2517] = 8'b11111111;
assign hamming[2518] = 8'b11111111;
assign hamming[2519] = 8'b11111111;
assign hamming[2520] = 8'b11011010;
assign hamming[2521] = 8'b10111010;
assign hamming[2522] = 8'b10001010;
assign hamming[2523] = 8'b10011010;
assign hamming[2524] = 8'b10011011;
assign hamming[2525] = 8'b10001011;
assign hamming[2526] = 8'b10111011;
assign hamming[2527] = 8'b11011011;
assign hamming[2528] = 8'b00011100;
assign hamming[2529] = 8'b11111111;
assign hamming[2530] = 8'b11111111;
assign hamming[2531] = 8'b11111111;
assign hamming[2532] = 8'b11111111;
assign hamming[2533] = 8'b11111111;
assign hamming[2534] = 8'b11111111;
assign hamming[2535] = 8'b00011101;
assign hamming[2536] = 8'b10011100;
assign hamming[2537] = 8'b10001100;
assign hamming[2538] = 8'b10111100;
assign hamming[2539] = 8'b11011100;
assign hamming[2540] = 8'b11011101;
assign hamming[2541] = 8'b10111101;
assign hamming[2542] = 8'b10001101;
assign hamming[2543] = 8'b10011101;
assign hamming[2544] = 8'b10001110;
assign hamming[2545] = 8'b10011110;
assign hamming[2546] = 8'b11011110;
assign hamming[2547] = 8'b10111110;
assign hamming[2548] = 8'b10111111;
assign hamming[2549] = 8'b11011111;
assign hamming[2550] = 8'b10011111;
assign hamming[2551] = 8'b10001111;
assign hamming[2552] = 8'b11111111;
assign hamming[2553] = 8'b00011110;
assign hamming[2554] = 8'b11111111;
assign hamming[2555] = 8'b11111111;
assign hamming[2556] = 8'b11111111;
assign hamming[2557] = 8'b11111111;
assign hamming[2558] = 8'b00011111;
assign hamming[2559] = 8'b11111111;
assign hamming[2560] = 8'b10100100;
assign hamming[2561] = 8'b10101000;
assign hamming[2562] = 8'b10100000;
assign hamming[2563] = 8'b10100010;
assign hamming[2564] = 8'b10100011;
assign hamming[2565] = 8'b10100001;
assign hamming[2566] = 8'b10101001;
assign hamming[2567] = 8'b10100101;
assign hamming[2568] = 8'b10100000;
assign hamming[2569] = 8'b10100001;
assign hamming[2570] = 8'b10100000;
assign hamming[2571] = 8'b10100000;
assign hamming[2572] = 8'b10100001;
assign hamming[2573] = 8'b10100001;
assign hamming[2574] = 8'b10100000;
assign hamming[2575] = 8'b10100001;
assign hamming[2576] = 8'b10100011;
assign hamming[2577] = 8'b10100010;
assign hamming[2578] = 8'b10100010;
assign hamming[2579] = 8'b10100010;
assign hamming[2580] = 8'b10100011;
assign hamming[2581] = 8'b10100011;
assign hamming[2582] = 8'b10100011;
assign hamming[2583] = 8'b10100010;
assign hamming[2584] = 8'b10101010;
assign hamming[2585] = 8'b10100110;
assign hamming[2586] = 8'b10100000;
assign hamming[2587] = 8'b10100010;
assign hamming[2588] = 8'b10100011;
assign hamming[2589] = 8'b10100001;
assign hamming[2590] = 8'b10100111;
assign hamming[2591] = 8'b10101011;
assign hamming[2592] = 8'b10100100;
assign hamming[2593] = 8'b10100100;
assign hamming[2594] = 8'b10100100;
assign hamming[2595] = 8'b10100101;
assign hamming[2596] = 8'b10100100;
assign hamming[2597] = 8'b10100101;
assign hamming[2598] = 8'b10100101;
assign hamming[2599] = 8'b10100101;
assign hamming[2600] = 8'b10100100;
assign hamming[2601] = 8'b10100110;
assign hamming[2602] = 8'b10100000;
assign hamming[2603] = 8'b10101100;
assign hamming[2604] = 8'b10101101;
assign hamming[2605] = 8'b10100001;
assign hamming[2606] = 8'b10100111;
assign hamming[2607] = 8'b10100101;
assign hamming[2608] = 8'b10100100;
assign hamming[2609] = 8'b10100110;
assign hamming[2610] = 8'b10101110;
assign hamming[2611] = 8'b10100010;
assign hamming[2612] = 8'b10100011;
assign hamming[2613] = 8'b10101111;
assign hamming[2614] = 8'b10100111;
assign hamming[2615] = 8'b10100101;
assign hamming[2616] = 8'b10100110;
assign hamming[2617] = 8'b10100110;
assign hamming[2618] = 8'b10100111;
assign hamming[2619] = 8'b10100110;
assign hamming[2620] = 8'b10100111;
assign hamming[2621] = 8'b10100110;
assign hamming[2622] = 8'b10100111;
assign hamming[2623] = 8'b10100111;
assign hamming[2624] = 8'b10101000;
assign hamming[2625] = 8'b10101000;
assign hamming[2626] = 8'b10101001;
assign hamming[2627] = 8'b10101000;
assign hamming[2628] = 8'b10101001;
assign hamming[2629] = 8'b10101000;
assign hamming[2630] = 8'b10101001;
assign hamming[2631] = 8'b10101001;
assign hamming[2632] = 8'b10101010;
assign hamming[2633] = 8'b10101000;
assign hamming[2634] = 8'b10100000;
assign hamming[2635] = 8'b10101100;
assign hamming[2636] = 8'b10101101;
assign hamming[2637] = 8'b10100001;
assign hamming[2638] = 8'b10101001;
assign hamming[2639] = 8'b10101011;
assign hamming[2640] = 8'b10101010;
assign hamming[2641] = 8'b10101000;
assign hamming[2642] = 8'b10101110;
assign hamming[2643] = 8'b10100010;
assign hamming[2644] = 8'b10100011;
assign hamming[2645] = 8'b10101111;
assign hamming[2646] = 8'b10101001;
assign hamming[2647] = 8'b10101011;
assign hamming[2648] = 8'b10101010;
assign hamming[2649] = 8'b10101010;
assign hamming[2650] = 8'b10101010;
assign hamming[2651] = 8'b10101011;
assign hamming[2652] = 8'b10101010;
assign hamming[2653] = 8'b10101011;
assign hamming[2654] = 8'b10101011;
assign hamming[2655] = 8'b10101011;
assign hamming[2656] = 8'b10100100;
assign hamming[2657] = 8'b10101000;
assign hamming[2658] = 8'b10101110;
assign hamming[2659] = 8'b10101100;
assign hamming[2660] = 8'b10101101;
assign hamming[2661] = 8'b10101111;
assign hamming[2662] = 8'b10101001;
assign hamming[2663] = 8'b10100101;
assign hamming[2664] = 8'b10101101;
assign hamming[2665] = 8'b10101100;
assign hamming[2666] = 8'b10101100;
assign hamming[2667] = 8'b10101100;
assign hamming[2668] = 8'b10101101;
assign hamming[2669] = 8'b10101101;
assign hamming[2670] = 8'b10101101;
assign hamming[2671] = 8'b10101100;
assign hamming[2672] = 8'b10101110;
assign hamming[2673] = 8'b10101111;
assign hamming[2674] = 8'b10101110;
assign hamming[2675] = 8'b10101110;
assign hamming[2676] = 8'b10101111;
assign hamming[2677] = 8'b10101111;
assign hamming[2678] = 8'b10101110;
assign hamming[2679] = 8'b10101111;
assign hamming[2680] = 8'b10101010;
assign hamming[2681] = 8'b10100110;
assign hamming[2682] = 8'b10101110;
assign hamming[2683] = 8'b10101100;
assign hamming[2684] = 8'b10101101;
assign hamming[2685] = 8'b10101111;
assign hamming[2686] = 8'b10100111;
assign hamming[2687] = 8'b10101011;
assign hamming[2688] = 8'b11111111;
assign hamming[2689] = 8'b11111111;
assign hamming[2690] = 8'b00100000;
assign hamming[2691] = 8'b11111111;
assign hamming[2692] = 8'b11111111;
assign hamming[2693] = 8'b00100001;
assign hamming[2694] = 8'b11111111;
assign hamming[2695] = 8'b11111111;
assign hamming[2696] = 8'b10000000;
assign hamming[2697] = 8'b11100000;
assign hamming[2698] = 8'b10100000;
assign hamming[2699] = 8'b10110000;
assign hamming[2700] = 8'b10110001;
assign hamming[2701] = 8'b10100001;
assign hamming[2702] = 8'b11100001;
assign hamming[2703] = 8'b10000001;
assign hamming[2704] = 8'b11100010;
assign hamming[2705] = 8'b10000010;
assign hamming[2706] = 8'b10110010;
assign hamming[2707] = 8'b10100010;
assign hamming[2708] = 8'b10100011;
assign hamming[2709] = 8'b10110011;
assign hamming[2710] = 8'b10000011;
assign hamming[2711] = 8'b11100011;
assign hamming[2712] = 8'b11111111;
assign hamming[2713] = 8'b11111111;
assign hamming[2714] = 8'b11111111;
assign hamming[2715] = 8'b00100010;
assign hamming[2716] = 8'b00100011;
assign hamming[2717] = 8'b11111111;
assign hamming[2718] = 8'b11111111;
assign hamming[2719] = 8'b11111111;
assign hamming[2720] = 8'b10100100;
assign hamming[2721] = 8'b10110100;
assign hamming[2722] = 8'b10000100;
assign hamming[2723] = 8'b11100100;
assign hamming[2724] = 8'b11100101;
assign hamming[2725] = 8'b10000101;
assign hamming[2726] = 8'b10110101;
assign hamming[2727] = 8'b10100101;
assign hamming[2728] = 8'b00100100;
assign hamming[2729] = 8'b11111111;
assign hamming[2730] = 8'b11111111;
assign hamming[2731] = 8'b11111111;
assign hamming[2732] = 8'b11111111;
assign hamming[2733] = 8'b11111111;
assign hamming[2734] = 8'b11111111;
assign hamming[2735] = 8'b00100101;
assign hamming[2736] = 8'b11111111;
assign hamming[2737] = 8'b00100110;
assign hamming[2738] = 8'b11111111;
assign hamming[2739] = 8'b11111111;
assign hamming[2740] = 8'b11111111;
assign hamming[2741] = 8'b11111111;
assign hamming[2742] = 8'b00100111;
assign hamming[2743] = 8'b11111111;
assign hamming[2744] = 8'b10110110;
assign hamming[2745] = 8'b10100110;
assign hamming[2746] = 8'b11100110;
assign hamming[2747] = 8'b10000110;
assign hamming[2748] = 8'b10000111;
assign hamming[2749] = 8'b11100111;
assign hamming[2750] = 8'b10100111;
assign hamming[2751] = 8'b10110111;
assign hamming[2752] = 8'b10111000;
assign hamming[2753] = 8'b10101000;
assign hamming[2754] = 8'b11101000;
assign hamming[2755] = 8'b10001000;
assign hamming[2756] = 8'b10001001;
assign hamming[2757] = 8'b11101001;
assign hamming[2758] = 8'b10101001;
assign hamming[2759] = 8'b10111001;
assign hamming[2760] = 8'b11111111;
assign hamming[2761] = 8'b00101000;
assign hamming[2762] = 8'b11111111;
assign hamming[2763] = 8'b11111111;
assign hamming[2764] = 8'b11111111;
assign hamming[2765] = 8'b11111111;
assign hamming[2766] = 8'b00101001;
assign hamming[2767] = 8'b11111111;
assign hamming[2768] = 8'b00101010;
assign hamming[2769] = 8'b11111111;
assign hamming[2770] = 8'b11111111;
assign hamming[2771] = 8'b11111111;
assign hamming[2772] = 8'b11111111;
assign hamming[2773] = 8'b11111111;
assign hamming[2774] = 8'b11111111;
assign hamming[2775] = 8'b00101011;
assign hamming[2776] = 8'b10101010;
assign hamming[2777] = 8'b10111010;
assign hamming[2778] = 8'b10001010;
assign hamming[2779] = 8'b11101010;
assign hamming[2780] = 8'b11101011;
assign hamming[2781] = 8'b10001011;
assign hamming[2782] = 8'b10111011;
assign hamming[2783] = 8'b10101011;
assign hamming[2784] = 8'b11111111;
assign hamming[2785] = 8'b11111111;
assign hamming[2786] = 8'b11111111;
assign hamming[2787] = 8'b00101100;
assign hamming[2788] = 8'b00101101;
assign hamming[2789] = 8'b11111111;
assign hamming[2790] = 8'b11111111;
assign hamming[2791] = 8'b11111111;
assign hamming[2792] = 8'b11101100;
assign hamming[2793] = 8'b10001100;
assign hamming[2794] = 8'b10111100;
assign hamming[2795] = 8'b10101100;
assign hamming[2796] = 8'b10101101;
assign hamming[2797] = 8'b10111101;
assign hamming[2798] = 8'b10001101;
assign hamming[2799] = 8'b11101101;
assign hamming[2800] = 8'b10001110;
assign hamming[2801] = 8'b11101110;
assign hamming[2802] = 8'b10101110;
assign hamming[2803] = 8'b10111110;
assign hamming[2804] = 8'b10111111;
assign hamming[2805] = 8'b10101111;
assign hamming[2806] = 8'b11101111;
assign hamming[2807] = 8'b10001111;
assign hamming[2808] = 8'b11111111;
assign hamming[2809] = 8'b11111111;
assign hamming[2810] = 8'b00101110;
assign hamming[2811] = 8'b11111111;
assign hamming[2812] = 8'b11111111;
assign hamming[2813] = 8'b00101111;
assign hamming[2814] = 8'b11111111;
assign hamming[2815] = 8'b11111111;
assign hamming[2816] = 8'b11111111;
assign hamming[2817] = 8'b11111111;
assign hamming[2818] = 8'b11111111;
assign hamming[2819] = 8'b00110000;
assign hamming[2820] = 8'b00110001;
assign hamming[2821] = 8'b11111111;
assign hamming[2822] = 8'b11111111;
assign hamming[2823] = 8'b11111111;
assign hamming[2824] = 8'b11110000;
assign hamming[2825] = 8'b10010000;
assign hamming[2826] = 8'b10100000;
assign hamming[2827] = 8'b10110000;
assign hamming[2828] = 8'b10110001;
assign hamming[2829] = 8'b10100001;
assign hamming[2830] = 8'b10010001;
assign hamming[2831] = 8'b11110001;
assign hamming[2832] = 8'b10010010;
assign hamming[2833] = 8'b11110010;
assign hamming[2834] = 8'b10110010;
assign hamming[2835] = 8'b10100010;
assign hamming[2836] = 8'b10100011;
assign hamming[2837] = 8'b10110011;
assign hamming[2838] = 8'b11110011;
assign hamming[2839] = 8'b10010011;
assign hamming[2840] = 8'b11111111;
assign hamming[2841] = 8'b11111111;
assign hamming[2842] = 8'b00110010;
assign hamming[2843] = 8'b11111111;
assign hamming[2844] = 8'b11111111;
assign hamming[2845] = 8'b00110011;
assign hamming[2846] = 8'b11111111;
assign hamming[2847] = 8'b11111111;
assign hamming[2848] = 8'b10100100;
assign hamming[2849] = 8'b10110100;
assign hamming[2850] = 8'b11110100;
assign hamming[2851] = 8'b10010100;
assign hamming[2852] = 8'b10010101;
assign hamming[2853] = 8'b11110101;
assign hamming[2854] = 8'b10110101;
assign hamming[2855] = 8'b10100101;
assign hamming[2856] = 8'b11111111;
assign hamming[2857] = 8'b00110100;
assign hamming[2858] = 8'b11111111;
assign hamming[2859] = 8'b11111111;
assign hamming[2860] = 8'b11111111;
assign hamming[2861] = 8'b11111111;
assign hamming[2862] = 8'b00110101;
assign hamming[2863] = 8'b11111111;
assign hamming[2864] = 8'b00110110;
assign hamming[2865] = 8'b11111111;
assign hamming[2866] = 8'b11111111;
assign hamming[2867] = 8'b11111111;
assign hamming[2868] = 8'b11111111;
assign hamming[2869] = 8'b11111111;
assign hamming[2870] = 8'b11111111;
assign hamming[2871] = 8'b00110111;
assign hamming[2872] = 8'b10110110;
assign hamming[2873] = 8'b10100110;
assign hamming[2874] = 8'b10010110;
assign hamming[2875] = 8'b11110110;
assign hamming[2876] = 8'b11110111;
assign hamming[2877] = 8'b10010111;
assign hamming[2878] = 8'b10100111;
assign hamming[2879] = 8'b10110111;
assign hamming[2880] = 8'b10111000;
assign hamming[2881] = 8'b10101000;
assign hamming[2882] = 8'b10011000;
assign hamming[2883] = 8'b11111000;
assign hamming[2884] = 8'b11111001;
assign hamming[2885] = 8'b10011001;
assign hamming[2886] = 8'b10101001;
assign hamming[2887] = 8'b10111001;
assign hamming[2888] = 8'b00111000;
assign hamming[2889] = 8'b11111111;
assign hamming[2890] = 8'b11111111;
assign hamming[2891] = 8'b11111111;
assign hamming[2892] = 8'b11111111;
assign hamming[2893] = 8'b11111111;
assign hamming[2894] = 8'b11111111;
assign hamming[2895] = 8'b00111001;
assign hamming[2896] = 8'b11111111;
assign hamming[2897] = 8'b00111010;
assign hamming[2898] = 8'b11111111;
assign hamming[2899] = 8'b11111111;
assign hamming[2900] = 8'b11111111;
assign hamming[2901] = 8'b11111111;
assign hamming[2902] = 8'b00111011;
assign hamming[2903] = 8'b11111111;
assign hamming[2904] = 8'b10101010;
assign hamming[2905] = 8'b10111010;
assign hamming[2906] = 8'b11111010;
assign hamming[2907] = 8'b10011010;
assign hamming[2908] = 8'b10011011;
assign hamming[2909] = 8'b11111011;
assign hamming[2910] = 8'b10111011;
assign hamming[2911] = 8'b10101011;
assign hamming[2912] = 8'b11111111;
assign hamming[2913] = 8'b11111111;
assign hamming[2914] = 8'b00111100;
assign hamming[2915] = 8'b11111111;
assign hamming[2916] = 8'b11111111;
assign hamming[2917] = 8'b00111101;
assign hamming[2918] = 8'b11111111;
assign hamming[2919] = 8'b11111111;
assign hamming[2920] = 8'b10011100;
assign hamming[2921] = 8'b11111100;
assign hamming[2922] = 8'b10111100;
assign hamming[2923] = 8'b10101100;
assign hamming[2924] = 8'b10101101;
assign hamming[2925] = 8'b10111101;
assign hamming[2926] = 8'b11111101;
assign hamming[2927] = 8'b10011101;
assign hamming[2928] = 8'b11111110;
assign hamming[2929] = 8'b10011110;
assign hamming[2930] = 8'b10101110;
assign hamming[2931] = 8'b10111110;
assign hamming[2932] = 8'b10111111;
assign hamming[2933] = 8'b10101111;
assign hamming[2934] = 8'b10011111;
assign hamming[2935] = 8'b11111111;
assign hamming[2936] = 8'b11111111;
assign hamming[2937] = 8'b11111111;
assign hamming[2938] = 8'b11111111;
assign hamming[2939] = 8'b00111110;
assign hamming[2940] = 8'b00111111;
assign hamming[2941] = 8'b11111111;
assign hamming[2942] = 8'b11111111;
assign hamming[2943] = 8'b11111111;
assign hamming[2944] = 8'b10111000;
assign hamming[2945] = 8'b10110100;
assign hamming[2946] = 8'b10110010;
assign hamming[2947] = 8'b10110000;
assign hamming[2948] = 8'b10110001;
assign hamming[2949] = 8'b10110011;
assign hamming[2950] = 8'b10110101;
assign hamming[2951] = 8'b10111001;
assign hamming[2952] = 8'b10110001;
assign hamming[2953] = 8'b10110000;
assign hamming[2954] = 8'b10110000;
assign hamming[2955] = 8'b10110000;
assign hamming[2956] = 8'b10110001;
assign hamming[2957] = 8'b10110001;
assign hamming[2958] = 8'b10110001;
assign hamming[2959] = 8'b10110000;
assign hamming[2960] = 8'b10110010;
assign hamming[2961] = 8'b10110011;
assign hamming[2962] = 8'b10110010;
assign hamming[2963] = 8'b10110010;
assign hamming[2964] = 8'b10110011;
assign hamming[2965] = 8'b10110011;
assign hamming[2966] = 8'b10110010;
assign hamming[2967] = 8'b10110011;
assign hamming[2968] = 8'b10110110;
assign hamming[2969] = 8'b10111010;
assign hamming[2970] = 8'b10110010;
assign hamming[2971] = 8'b10110000;
assign hamming[2972] = 8'b10110001;
assign hamming[2973] = 8'b10110011;
assign hamming[2974] = 8'b10111011;
assign hamming[2975] = 8'b10110111;
assign hamming[2976] = 8'b10110100;
assign hamming[2977] = 8'b10110100;
assign hamming[2978] = 8'b10110101;
assign hamming[2979] = 8'b10110100;
assign hamming[2980] = 8'b10110101;
assign hamming[2981] = 8'b10110100;
assign hamming[2982] = 8'b10110101;
assign hamming[2983] = 8'b10110101;
assign hamming[2984] = 8'b10110110;
assign hamming[2985] = 8'b10110100;
assign hamming[2986] = 8'b10111100;
assign hamming[2987] = 8'b10110000;
assign hamming[2988] = 8'b10110001;
assign hamming[2989] = 8'b10111101;
assign hamming[2990] = 8'b10110101;
assign hamming[2991] = 8'b10110111;
assign hamming[2992] = 8'b10110110;
assign hamming[2993] = 8'b10110100;
assign hamming[2994] = 8'b10110010;
assign hamming[2995] = 8'b10111110;
assign hamming[2996] = 8'b10111111;
assign hamming[2997] = 8'b10110011;
assign hamming[2998] = 8'b10110101;
assign hamming[2999] = 8'b10110111;
assign hamming[3000] = 8'b10110110;
assign hamming[3001] = 8'b10110110;
assign hamming[3002] = 8'b10110110;
assign hamming[3003] = 8'b10110111;
assign hamming[3004] = 8'b10110110;
assign hamming[3005] = 8'b10110111;
assign hamming[3006] = 8'b10110111;
assign hamming[3007] = 8'b10110111;
assign hamming[3008] = 8'b10111000;
assign hamming[3009] = 8'b10111000;
assign hamming[3010] = 8'b10111000;
assign hamming[3011] = 8'b10111001;
assign hamming[3012] = 8'b10111000;
assign hamming[3013] = 8'b10111001;
assign hamming[3014] = 8'b10111001;
assign hamming[3015] = 8'b10111001;
assign hamming[3016] = 8'b10111000;
assign hamming[3017] = 8'b10111010;
assign hamming[3018] = 8'b10111100;
assign hamming[3019] = 8'b10110000;
assign hamming[3020] = 8'b10110001;
assign hamming[3021] = 8'b10111101;
assign hamming[3022] = 8'b10111011;
assign hamming[3023] = 8'b10111001;
assign hamming[3024] = 8'b10111000;
assign hamming[3025] = 8'b10111010;
assign hamming[3026] = 8'b10110010;
assign hamming[3027] = 8'b10111110;
assign hamming[3028] = 8'b10111111;
assign hamming[3029] = 8'b10110011;
assign hamming[3030] = 8'b10111011;
assign hamming[3031] = 8'b10111001;
assign hamming[3032] = 8'b10111010;
assign hamming[3033] = 8'b10111010;
assign hamming[3034] = 8'b10111011;
assign hamming[3035] = 8'b10111010;
assign hamming[3036] = 8'b10111011;
assign hamming[3037] = 8'b10111010;
assign hamming[3038] = 8'b10111011;
assign hamming[3039] = 8'b10111011;
assign hamming[3040] = 8'b10111000;
assign hamming[3041] = 8'b10110100;
assign hamming[3042] = 8'b10111100;
assign hamming[3043] = 8'b10111110;
assign hamming[3044] = 8'b10111111;
assign hamming[3045] = 8'b10111101;
assign hamming[3046] = 8'b10110101;
assign hamming[3047] = 8'b10111001;
assign hamming[3048] = 8'b10111100;
assign hamming[3049] = 8'b10111101;
assign hamming[3050] = 8'b10111100;
assign hamming[3051] = 8'b10111100;
assign hamming[3052] = 8'b10111101;
assign hamming[3053] = 8'b10111101;
assign hamming[3054] = 8'b10111100;
assign hamming[3055] = 8'b10111101;
assign hamming[3056] = 8'b10111111;
assign hamming[3057] = 8'b10111110;
assign hamming[3058] = 8'b10111110;
assign hamming[3059] = 8'b10111110;
assign hamming[3060] = 8'b10111111;
assign hamming[3061] = 8'b10111111;
assign hamming[3062] = 8'b10111111;
assign hamming[3063] = 8'b10111110;
assign hamming[3064] = 8'b10110110;
assign hamming[3065] = 8'b10111010;
assign hamming[3066] = 8'b10111100;
assign hamming[3067] = 8'b10111110;
assign hamming[3068] = 8'b10111111;
assign hamming[3069] = 8'b10111101;
assign hamming[3070] = 8'b10111011;
assign hamming[3071] = 8'b10110111;
assign hamming[3072] = 8'b11001000;
assign hamming[3073] = 8'b11000100;
assign hamming[3074] = 8'b11000010;
assign hamming[3075] = 8'b11000000;
assign hamming[3076] = 8'b11000001;
assign hamming[3077] = 8'b11000011;
assign hamming[3078] = 8'b11000101;
assign hamming[3079] = 8'b11001001;
assign hamming[3080] = 8'b11000001;
assign hamming[3081] = 8'b11000000;
assign hamming[3082] = 8'b11000000;
assign hamming[3083] = 8'b11000000;
assign hamming[3084] = 8'b11000001;
assign hamming[3085] = 8'b11000001;
assign hamming[3086] = 8'b11000001;
assign hamming[3087] = 8'b11000000;
assign hamming[3088] = 8'b11000010;
assign hamming[3089] = 8'b11000011;
assign hamming[3090] = 8'b11000010;
assign hamming[3091] = 8'b11000010;
assign hamming[3092] = 8'b11000011;
assign hamming[3093] = 8'b11000011;
assign hamming[3094] = 8'b11000010;
assign hamming[3095] = 8'b11000011;
assign hamming[3096] = 8'b11000110;
assign hamming[3097] = 8'b11001010;
assign hamming[3098] = 8'b11000010;
assign hamming[3099] = 8'b11000000;
assign hamming[3100] = 8'b11000001;
assign hamming[3101] = 8'b11000011;
assign hamming[3102] = 8'b11001011;
assign hamming[3103] = 8'b11000111;
assign hamming[3104] = 8'b11000100;
assign hamming[3105] = 8'b11000100;
assign hamming[3106] = 8'b11000101;
assign hamming[3107] = 8'b11000100;
assign hamming[3108] = 8'b11000101;
assign hamming[3109] = 8'b11000100;
assign hamming[3110] = 8'b11000101;
assign hamming[3111] = 8'b11000101;
assign hamming[3112] = 8'b11000110;
assign hamming[3113] = 8'b11000100;
assign hamming[3114] = 8'b11001100;
assign hamming[3115] = 8'b11000000;
assign hamming[3116] = 8'b11000001;
assign hamming[3117] = 8'b11001101;
assign hamming[3118] = 8'b11000101;
assign hamming[3119] = 8'b11000111;
assign hamming[3120] = 8'b11000110;
assign hamming[3121] = 8'b11000100;
assign hamming[3122] = 8'b11000010;
assign hamming[3123] = 8'b11001110;
assign hamming[3124] = 8'b11001111;
assign hamming[3125] = 8'b11000011;
assign hamming[3126] = 8'b11000101;
assign hamming[3127] = 8'b11000111;
assign hamming[3128] = 8'b11000110;
assign hamming[3129] = 8'b11000110;
assign hamming[3130] = 8'b11000110;
assign hamming[3131] = 8'b11000111;
assign hamming[3132] = 8'b11000110;
assign hamming[3133] = 8'b11000111;
assign hamming[3134] = 8'b11000111;
assign hamming[3135] = 8'b11000111;
assign hamming[3136] = 8'b11001000;
assign hamming[3137] = 8'b11001000;
assign hamming[3138] = 8'b11001000;
assign hamming[3139] = 8'b11001001;
assign hamming[3140] = 8'b11001000;
assign hamming[3141] = 8'b11001001;
assign hamming[3142] = 8'b11001001;
assign hamming[3143] = 8'b11001001;
assign hamming[3144] = 8'b11001000;
assign hamming[3145] = 8'b11001010;
assign hamming[3146] = 8'b11001100;
assign hamming[3147] = 8'b11000000;
assign hamming[3148] = 8'b11000001;
assign hamming[3149] = 8'b11001101;
assign hamming[3150] = 8'b11001011;
assign hamming[3151] = 8'b11001001;
assign hamming[3152] = 8'b11001000;
assign hamming[3153] = 8'b11001010;
assign hamming[3154] = 8'b11000010;
assign hamming[3155] = 8'b11001110;
assign hamming[3156] = 8'b11001111;
assign hamming[3157] = 8'b11000011;
assign hamming[3158] = 8'b11001011;
assign hamming[3159] = 8'b11001001;
assign hamming[3160] = 8'b11001010;
assign hamming[3161] = 8'b11001010;
assign hamming[3162] = 8'b11001011;
assign hamming[3163] = 8'b11001010;
assign hamming[3164] = 8'b11001011;
assign hamming[3165] = 8'b11001010;
assign hamming[3166] = 8'b11001011;
assign hamming[3167] = 8'b11001011;
assign hamming[3168] = 8'b11001000;
assign hamming[3169] = 8'b11000100;
assign hamming[3170] = 8'b11001100;
assign hamming[3171] = 8'b11001110;
assign hamming[3172] = 8'b11001111;
assign hamming[3173] = 8'b11001101;
assign hamming[3174] = 8'b11000101;
assign hamming[3175] = 8'b11001001;
assign hamming[3176] = 8'b11001100;
assign hamming[3177] = 8'b11001101;
assign hamming[3178] = 8'b11001100;
assign hamming[3179] = 8'b11001100;
assign hamming[3180] = 8'b11001101;
assign hamming[3181] = 8'b11001101;
assign hamming[3182] = 8'b11001100;
assign hamming[3183] = 8'b11001101;
assign hamming[3184] = 8'b11001111;
assign hamming[3185] = 8'b11001110;
assign hamming[3186] = 8'b11001110;
assign hamming[3187] = 8'b11001110;
assign hamming[3188] = 8'b11001111;
assign hamming[3189] = 8'b11001111;
assign hamming[3190] = 8'b11001111;
assign hamming[3191] = 8'b11001110;
assign hamming[3192] = 8'b11000110;
assign hamming[3193] = 8'b11001010;
assign hamming[3194] = 8'b11001100;
assign hamming[3195] = 8'b11001110;
assign hamming[3196] = 8'b11001111;
assign hamming[3197] = 8'b11001101;
assign hamming[3198] = 8'b11001011;
assign hamming[3199] = 8'b11000111;
assign hamming[3200] = 8'b11111111;
assign hamming[3201] = 8'b11111111;
assign hamming[3202] = 8'b11111111;
assign hamming[3203] = 8'b01000000;
assign hamming[3204] = 8'b01000001;
assign hamming[3205] = 8'b11111111;
assign hamming[3206] = 8'b11111111;
assign hamming[3207] = 8'b11111111;
assign hamming[3208] = 8'b10000000;
assign hamming[3209] = 8'b11100000;
assign hamming[3210] = 8'b11010000;
assign hamming[3211] = 8'b11000000;
assign hamming[3212] = 8'b11000001;
assign hamming[3213] = 8'b11010001;
assign hamming[3214] = 8'b11100001;
assign hamming[3215] = 8'b10000001;
assign hamming[3216] = 8'b11100010;
assign hamming[3217] = 8'b10000010;
assign hamming[3218] = 8'b11000010;
assign hamming[3219] = 8'b11010010;
assign hamming[3220] = 8'b11010011;
assign hamming[3221] = 8'b11000011;
assign hamming[3222] = 8'b10000011;
assign hamming[3223] = 8'b11100011;
assign hamming[3224] = 8'b11111111;
assign hamming[3225] = 8'b11111111;
assign hamming[3226] = 8'b01000010;
assign hamming[3227] = 8'b11111111;
assign hamming[3228] = 8'b11111111;
assign hamming[3229] = 8'b01000011;
assign hamming[3230] = 8'b11111111;
assign hamming[3231] = 8'b11111111;
assign hamming[3232] = 8'b11010100;
assign hamming[3233] = 8'b11000100;
assign hamming[3234] = 8'b10000100;
assign hamming[3235] = 8'b11100100;
assign hamming[3236] = 8'b11100101;
assign hamming[3237] = 8'b10000101;
assign hamming[3238] = 8'b11000101;
assign hamming[3239] = 8'b11010101;
assign hamming[3240] = 8'b11111111;
assign hamming[3241] = 8'b01000100;
assign hamming[3242] = 8'b11111111;
assign hamming[3243] = 8'b11111111;
assign hamming[3244] = 8'b11111111;
assign hamming[3245] = 8'b11111111;
assign hamming[3246] = 8'b01000101;
assign hamming[3247] = 8'b11111111;
assign hamming[3248] = 8'b01000110;
assign hamming[3249] = 8'b11111111;
assign hamming[3250] = 8'b11111111;
assign hamming[3251] = 8'b11111111;
assign hamming[3252] = 8'b11111111;
assign hamming[3253] = 8'b11111111;
assign hamming[3254] = 8'b11111111;
assign hamming[3255] = 8'b01000111;
assign hamming[3256] = 8'b11000110;
assign hamming[3257] = 8'b11010110;
assign hamming[3258] = 8'b11100110;
assign hamming[3259] = 8'b10000110;
assign hamming[3260] = 8'b10000111;
assign hamming[3261] = 8'b11100111;
assign hamming[3262] = 8'b11010111;
assign hamming[3263] = 8'b11000111;
assign hamming[3264] = 8'b11001000;
assign hamming[3265] = 8'b11011000;
assign hamming[3266] = 8'b11101000;
assign hamming[3267] = 8'b10001000;
assign hamming[3268] = 8'b10001001;
assign hamming[3269] = 8'b11101001;
assign hamming[3270] = 8'b11011001;
assign hamming[3271] = 8'b11001001;
assign hamming[3272] = 8'b01001000;
assign hamming[3273] = 8'b11111111;
assign hamming[3274] = 8'b11111111;
assign hamming[3275] = 8'b11111111;
assign hamming[3276] = 8'b11111111;
assign hamming[3277] = 8'b11111111;
assign hamming[3278] = 8'b11111111;
assign hamming[3279] = 8'b01001001;
assign hamming[3280] = 8'b11111111;
assign hamming[3281] = 8'b01001010;
assign hamming[3282] = 8'b11111111;
assign hamming[3283] = 8'b11111111;
assign hamming[3284] = 8'b11111111;
assign hamming[3285] = 8'b11111111;
assign hamming[3286] = 8'b01001011;
assign hamming[3287] = 8'b11111111;
assign hamming[3288] = 8'b11011010;
assign hamming[3289] = 8'b11001010;
assign hamming[3290] = 8'b10001010;
assign hamming[3291] = 8'b11101010;
assign hamming[3292] = 8'b11101011;
assign hamming[3293] = 8'b10001011;
assign hamming[3294] = 8'b11001011;
assign hamming[3295] = 8'b11011011;
assign hamming[3296] = 8'b11111111;
assign hamming[3297] = 8'b11111111;
assign hamming[3298] = 8'b01001100;
assign hamming[3299] = 8'b11111111;
assign hamming[3300] = 8'b11111111;
assign hamming[3301] = 8'b01001101;
assign hamming[3302] = 8'b11111111;
assign hamming[3303] = 8'b11111111;
assign hamming[3304] = 8'b11101100;
assign hamming[3305] = 8'b10001100;
assign hamming[3306] = 8'b11001100;
assign hamming[3307] = 8'b11011100;
assign hamming[3308] = 8'b11011101;
assign hamming[3309] = 8'b11001101;
assign hamming[3310] = 8'b10001101;
assign hamming[3311] = 8'b11101101;
assign hamming[3312] = 8'b10001110;
assign hamming[3313] = 8'b11101110;
assign hamming[3314] = 8'b11011110;
assign hamming[3315] = 8'b11001110;
assign hamming[3316] = 8'b11001111;
assign hamming[3317] = 8'b11011111;
assign hamming[3318] = 8'b11101111;
assign hamming[3319] = 8'b10001111;
assign hamming[3320] = 8'b11111111;
assign hamming[3321] = 8'b11111111;
assign hamming[3322] = 8'b11111111;
assign hamming[3323] = 8'b01001110;
assign hamming[3324] = 8'b01001111;
assign hamming[3325] = 8'b11111111;
assign hamming[3326] = 8'b11111111;
assign hamming[3327] = 8'b11111111;
assign hamming[3328] = 8'b11111111;
assign hamming[3329] = 8'b11111111;
assign hamming[3330] = 8'b01010000;
assign hamming[3331] = 8'b11111111;
assign hamming[3332] = 8'b11111111;
assign hamming[3333] = 8'b01010001;
assign hamming[3334] = 8'b11111111;
assign hamming[3335] = 8'b11111111;
assign hamming[3336] = 8'b11110000;
assign hamming[3337] = 8'b10010000;
assign hamming[3338] = 8'b11010000;
assign hamming[3339] = 8'b11000000;
assign hamming[3340] = 8'b11000001;
assign hamming[3341] = 8'b11010001;
assign hamming[3342] = 8'b10010001;
assign hamming[3343] = 8'b11110001;
assign hamming[3344] = 8'b10010010;
assign hamming[3345] = 8'b11110010;
assign hamming[3346] = 8'b11000010;
assign hamming[3347] = 8'b11010010;
assign hamming[3348] = 8'b11010011;
assign hamming[3349] = 8'b11000011;
assign hamming[3350] = 8'b11110011;
assign hamming[3351] = 8'b10010011;
assign hamming[3352] = 8'b11111111;
assign hamming[3353] = 8'b11111111;
assign hamming[3354] = 8'b11111111;
assign hamming[3355] = 8'b01010010;
assign hamming[3356] = 8'b01010011;
assign hamming[3357] = 8'b11111111;
assign hamming[3358] = 8'b11111111;
assign hamming[3359] = 8'b11111111;
assign hamming[3360] = 8'b11010100;
assign hamming[3361] = 8'b11000100;
assign hamming[3362] = 8'b11110100;
assign hamming[3363] = 8'b10010100;
assign hamming[3364] = 8'b10010101;
assign hamming[3365] = 8'b11110101;
assign hamming[3366] = 8'b11000101;
assign hamming[3367] = 8'b11010101;
assign hamming[3368] = 8'b01010100;
assign hamming[3369] = 8'b11111111;
assign hamming[3370] = 8'b11111111;
assign hamming[3371] = 8'b11111111;
assign hamming[3372] = 8'b11111111;
assign hamming[3373] = 8'b11111111;
assign hamming[3374] = 8'b11111111;
assign hamming[3375] = 8'b01010101;
assign hamming[3376] = 8'b11111111;
assign hamming[3377] = 8'b01010110;
assign hamming[3378] = 8'b11111111;
assign hamming[3379] = 8'b11111111;
assign hamming[3380] = 8'b11111111;
assign hamming[3381] = 8'b11111111;
assign hamming[3382] = 8'b01010111;
assign hamming[3383] = 8'b11111111;
assign hamming[3384] = 8'b11000110;
assign hamming[3385] = 8'b11010110;
assign hamming[3386] = 8'b10010110;
assign hamming[3387] = 8'b11110110;
assign hamming[3388] = 8'b11110111;
assign hamming[3389] = 8'b10010111;
assign hamming[3390] = 8'b11010111;
assign hamming[3391] = 8'b11000111;
assign hamming[3392] = 8'b11001000;
assign hamming[3393] = 8'b11011000;
assign hamming[3394] = 8'b10011000;
assign hamming[3395] = 8'b11111000;
assign hamming[3396] = 8'b11111001;
assign hamming[3397] = 8'b10011001;
assign hamming[3398] = 8'b11011001;
assign hamming[3399] = 8'b11001001;
assign hamming[3400] = 8'b11111111;
assign hamming[3401] = 8'b01011000;
assign hamming[3402] = 8'b11111111;
assign hamming[3403] = 8'b11111111;
assign hamming[3404] = 8'b11111111;
assign hamming[3405] = 8'b11111111;
assign hamming[3406] = 8'b01011001;
assign hamming[3407] = 8'b11111111;
assign hamming[3408] = 8'b01011010;
assign hamming[3409] = 8'b11111111;
assign hamming[3410] = 8'b11111111;
assign hamming[3411] = 8'b11111111;
assign hamming[3412] = 8'b11111111;
assign hamming[3413] = 8'b11111111;
assign hamming[3414] = 8'b11111111;
assign hamming[3415] = 8'b01011011;
assign hamming[3416] = 8'b11011010;
assign hamming[3417] = 8'b11001010;
assign hamming[3418] = 8'b11111010;
assign hamming[3419] = 8'b10011010;
assign hamming[3420] = 8'b10011011;
assign hamming[3421] = 8'b11111011;
assign hamming[3422] = 8'b11001011;
assign hamming[3423] = 8'b11011011;
assign hamming[3424] = 8'b11111111;
assign hamming[3425] = 8'b11111111;
assign hamming[3426] = 8'b11111111;
assign hamming[3427] = 8'b01011100;
assign hamming[3428] = 8'b01011101;
assign hamming[3429] = 8'b11111111;
assign hamming[3430] = 8'b11111111;
assign hamming[3431] = 8'b11111111;
assign hamming[3432] = 8'b10011100;
assign hamming[3433] = 8'b11111100;
assign hamming[3434] = 8'b11001100;
assign hamming[3435] = 8'b11011100;
assign hamming[3436] = 8'b11011101;
assign hamming[3437] = 8'b11001101;
assign hamming[3438] = 8'b11111101;
assign hamming[3439] = 8'b10011101;
assign hamming[3440] = 8'b11111110;
assign hamming[3441] = 8'b10011110;
assign hamming[3442] = 8'b11011110;
assign hamming[3443] = 8'b11001110;
assign hamming[3444] = 8'b11001111;
assign hamming[3445] = 8'b11011111;
assign hamming[3446] = 8'b10011111;
assign hamming[3447] = 8'b11111111;
assign hamming[3448] = 8'b11111111;
assign hamming[3449] = 8'b11111111;
assign hamming[3450] = 8'b01011110;
assign hamming[3451] = 8'b11111111;
assign hamming[3452] = 8'b11111111;
assign hamming[3453] = 8'b01011111;
assign hamming[3454] = 8'b11111111;
assign hamming[3455] = 8'b11111111;
assign hamming[3456] = 8'b11010100;
assign hamming[3457] = 8'b11011000;
assign hamming[3458] = 8'b11010000;
assign hamming[3459] = 8'b11010010;
assign hamming[3460] = 8'b11010011;
assign hamming[3461] = 8'b11010001;
assign hamming[3462] = 8'b11011001;
assign hamming[3463] = 8'b11010101;
assign hamming[3464] = 8'b11010000;
assign hamming[3465] = 8'b11010001;
assign hamming[3466] = 8'b11010000;
assign hamming[3467] = 8'b11010000;
assign hamming[3468] = 8'b11010001;
assign hamming[3469] = 8'b11010001;
assign hamming[3470] = 8'b11010000;
assign hamming[3471] = 8'b11010001;
assign hamming[3472] = 8'b11010011;
assign hamming[3473] = 8'b11010010;
assign hamming[3474] = 8'b11010010;
assign hamming[3475] = 8'b11010010;
assign hamming[3476] = 8'b11010011;
assign hamming[3477] = 8'b11010011;
assign hamming[3478] = 8'b11010011;
assign hamming[3479] = 8'b11010010;
assign hamming[3480] = 8'b11011010;
assign hamming[3481] = 8'b11010110;
assign hamming[3482] = 8'b11010000;
assign hamming[3483] = 8'b11010010;
assign hamming[3484] = 8'b11010011;
assign hamming[3485] = 8'b11010001;
assign hamming[3486] = 8'b11010111;
assign hamming[3487] = 8'b11011011;
assign hamming[3488] = 8'b11010100;
assign hamming[3489] = 8'b11010100;
assign hamming[3490] = 8'b11010100;
assign hamming[3491] = 8'b11010101;
assign hamming[3492] = 8'b11010100;
assign hamming[3493] = 8'b11010101;
assign hamming[3494] = 8'b11010101;
assign hamming[3495] = 8'b11010101;
assign hamming[3496] = 8'b11010100;
assign hamming[3497] = 8'b11010110;
assign hamming[3498] = 8'b11010000;
assign hamming[3499] = 8'b11011100;
assign hamming[3500] = 8'b11011101;
assign hamming[3501] = 8'b11010001;
assign hamming[3502] = 8'b11010111;
assign hamming[3503] = 8'b11010101;
assign hamming[3504] = 8'b11010100;
assign hamming[3505] = 8'b11010110;
assign hamming[3506] = 8'b11011110;
assign hamming[3507] = 8'b11010010;
assign hamming[3508] = 8'b11010011;
assign hamming[3509] = 8'b11011111;
assign hamming[3510] = 8'b11010111;
assign hamming[3511] = 8'b11010101;
assign hamming[3512] = 8'b11010110;
assign hamming[3513] = 8'b11010110;
assign hamming[3514] = 8'b11010111;
assign hamming[3515] = 8'b11010110;
assign hamming[3516] = 8'b11010111;
assign hamming[3517] = 8'b11010110;
assign hamming[3518] = 8'b11010111;
assign hamming[3519] = 8'b11010111;
assign hamming[3520] = 8'b11011000;
assign hamming[3521] = 8'b11011000;
assign hamming[3522] = 8'b11011001;
assign hamming[3523] = 8'b11011000;
assign hamming[3524] = 8'b11011001;
assign hamming[3525] = 8'b11011000;
assign hamming[3526] = 8'b11011001;
assign hamming[3527] = 8'b11011001;
assign hamming[3528] = 8'b11011010;
assign hamming[3529] = 8'b11011000;
assign hamming[3530] = 8'b11010000;
assign hamming[3531] = 8'b11011100;
assign hamming[3532] = 8'b11011101;
assign hamming[3533] = 8'b11010001;
assign hamming[3534] = 8'b11011001;
assign hamming[3535] = 8'b11011011;
assign hamming[3536] = 8'b11011010;
assign hamming[3537] = 8'b11011000;
assign hamming[3538] = 8'b11011110;
assign hamming[3539] = 8'b11010010;
assign hamming[3540] = 8'b11010011;
assign hamming[3541] = 8'b11011111;
assign hamming[3542] = 8'b11011001;
assign hamming[3543] = 8'b11011011;
assign hamming[3544] = 8'b11011010;
assign hamming[3545] = 8'b11011010;
assign hamming[3546] = 8'b11011010;
assign hamming[3547] = 8'b11011011;
assign hamming[3548] = 8'b11011010;
assign hamming[3549] = 8'b11011011;
assign hamming[3550] = 8'b11011011;
assign hamming[3551] = 8'b11011011;
assign hamming[3552] = 8'b11010100;
assign hamming[3553] = 8'b11011000;
assign hamming[3554] = 8'b11011110;
assign hamming[3555] = 8'b11011100;
assign hamming[3556] = 8'b11011101;
assign hamming[3557] = 8'b11011111;
assign hamming[3558] = 8'b11011001;
assign hamming[3559] = 8'b11010101;
assign hamming[3560] = 8'b11011101;
assign hamming[3561] = 8'b11011100;
assign hamming[3562] = 8'b11011100;
assign hamming[3563] = 8'b11011100;
assign hamming[3564] = 8'b11011101;
assign hamming[3565] = 8'b11011101;
assign hamming[3566] = 8'b11011101;
assign hamming[3567] = 8'b11011100;
assign hamming[3568] = 8'b11011110;
assign hamming[3569] = 8'b11011111;
assign hamming[3570] = 8'b11011110;
assign hamming[3571] = 8'b11011110;
assign hamming[3572] = 8'b11011111;
assign hamming[3573] = 8'b11011111;
assign hamming[3574] = 8'b11011110;
assign hamming[3575] = 8'b11011111;
assign hamming[3576] = 8'b11011010;
assign hamming[3577] = 8'b11010110;
assign hamming[3578] = 8'b11011110;
assign hamming[3579] = 8'b11011100;
assign hamming[3580] = 8'b11011101;
assign hamming[3581] = 8'b11011111;
assign hamming[3582] = 8'b11010111;
assign hamming[3583] = 8'b11011011;
assign hamming[3584] = 8'b11111111;
assign hamming[3585] = 8'b01100000;
assign hamming[3586] = 8'b11111111;
assign hamming[3587] = 8'b11111111;
assign hamming[3588] = 8'b11111111;
assign hamming[3589] = 8'b11111111;
assign hamming[3590] = 8'b01100001;
assign hamming[3591] = 8'b11111111;
assign hamming[3592] = 8'b11110000;
assign hamming[3593] = 8'b11100000;
assign hamming[3594] = 8'b10100000;
assign hamming[3595] = 8'b11000000;
assign hamming[3596] = 8'b11000001;
assign hamming[3597] = 8'b10100001;
assign hamming[3598] = 8'b11100001;
assign hamming[3599] = 8'b11110001;
assign hamming[3600] = 8'b11100010;
assign hamming[3601] = 8'b11110010;
assign hamming[3602] = 8'b11000010;
assign hamming[3603] = 8'b10100010;
assign hamming[3604] = 8'b10100011;
assign hamming[3605] = 8'b11000011;
assign hamming[3606] = 8'b11110011;
assign hamming[3607] = 8'b11100011;
assign hamming[3608] = 8'b01100010;
assign hamming[3609] = 8'b11111111;
assign hamming[3610] = 8'b11111111;
assign hamming[3611] = 8'b11111111;
assign hamming[3612] = 8'b11111111;
assign hamming[3613] = 8'b11111111;
assign hamming[3614] = 8'b11111111;
assign hamming[3615] = 8'b01100011;
assign hamming[3616] = 8'b10100100;
assign hamming[3617] = 8'b11000100;
assign hamming[3618] = 8'b11110100;
assign hamming[3619] = 8'b11100100;
assign hamming[3620] = 8'b11100101;
assign hamming[3621] = 8'b11110101;
assign hamming[3622] = 8'b11000101;
assign hamming[3623] = 8'b10100101;
assign hamming[3624] = 8'b11111111;
assign hamming[3625] = 8'b11111111;
assign hamming[3626] = 8'b11111111;
assign hamming[3627] = 8'b01100100;
assign hamming[3628] = 8'b01100101;
assign hamming[3629] = 8'b11111111;
assign hamming[3630] = 8'b11111111;
assign hamming[3631] = 8'b11111111;
assign hamming[3632] = 8'b11111111;
assign hamming[3633] = 8'b11111111;
assign hamming[3634] = 8'b01100110;
assign hamming[3635] = 8'b11111111;
assign hamming[3636] = 8'b11111111;
assign hamming[3637] = 8'b01100111;
assign hamming[3638] = 8'b11111111;
assign hamming[3639] = 8'b11111111;
assign hamming[3640] = 8'b11000110;
assign hamming[3641] = 8'b10100110;
assign hamming[3642] = 8'b11100110;
assign hamming[3643] = 8'b11110110;
assign hamming[3644] = 8'b11110111;
assign hamming[3645] = 8'b11100111;
assign hamming[3646] = 8'b10100111;
assign hamming[3647] = 8'b11000111;
assign hamming[3648] = 8'b11001000;
assign hamming[3649] = 8'b10101000;
assign hamming[3650] = 8'b11101000;
assign hamming[3651] = 8'b11111000;
assign hamming[3652] = 8'b11111001;
assign hamming[3653] = 8'b11101001;
assign hamming[3654] = 8'b10101001;
assign hamming[3655] = 8'b11001001;
assign hamming[3656] = 8'b11111111;
assign hamming[3657] = 8'b11111111;
assign hamming[3658] = 8'b01101000;
assign hamming[3659] = 8'b11111111;
assign hamming[3660] = 8'b11111111;
assign hamming[3661] = 8'b01101001;
assign hamming[3662] = 8'b11111111;
assign hamming[3663] = 8'b11111111;
assign hamming[3664] = 8'b11111111;
assign hamming[3665] = 8'b11111111;
assign hamming[3666] = 8'b11111111;
assign hamming[3667] = 8'b01101010;
assign hamming[3668] = 8'b01101011;
assign hamming[3669] = 8'b11111111;
assign hamming[3670] = 8'b11111111;
assign hamming[3671] = 8'b11111111;
assign hamming[3672] = 8'b10101010;
assign hamming[3673] = 8'b11001010;
assign hamming[3674] = 8'b11111010;
assign hamming[3675] = 8'b11101010;
assign hamming[3676] = 8'b11101011;
assign hamming[3677] = 8'b11111011;
assign hamming[3678] = 8'b11001011;
assign hamming[3679] = 8'b10101011;
assign hamming[3680] = 8'b01101100;
assign hamming[3681] = 8'b11111111;
assign hamming[3682] = 8'b11111111;
assign hamming[3683] = 8'b11111111;
assign hamming[3684] = 8'b11111111;
assign hamming[3685] = 8'b11111111;
assign hamming[3686] = 8'b11111111;
assign hamming[3687] = 8'b01101101;
assign hamming[3688] = 8'b11101100;
assign hamming[3689] = 8'b11111100;
assign hamming[3690] = 8'b11001100;
assign hamming[3691] = 8'b10101100;
assign hamming[3692] = 8'b10101101;
assign hamming[3693] = 8'b11001101;
assign hamming[3694] = 8'b11111101;
assign hamming[3695] = 8'b11101101;
assign hamming[3696] = 8'b11111110;
assign hamming[3697] = 8'b11101110;
assign hamming[3698] = 8'b10101110;
assign hamming[3699] = 8'b11001110;
assign hamming[3700] = 8'b11001111;
assign hamming[3701] = 8'b10101111;
assign hamming[3702] = 8'b11101111;
assign hamming[3703] = 8'b11111111;
assign hamming[3704] = 8'b11111111;
assign hamming[3705] = 8'b01101110;
assign hamming[3706] = 8'b11111111;
assign hamming[3707] = 8'b11111111;
assign hamming[3708] = 8'b11111111;
assign hamming[3709] = 8'b11111111;
assign hamming[3710] = 8'b01101111;
assign hamming[3711] = 8'b11111111;
assign hamming[3712] = 8'b11100010;
assign hamming[3713] = 8'b11100000;
assign hamming[3714] = 8'b11101000;
assign hamming[3715] = 8'b11100100;
assign hamming[3716] = 8'b11100101;
assign hamming[3717] = 8'b11101001;
assign hamming[3718] = 8'b11100001;
assign hamming[3719] = 8'b11100011;
assign hamming[3720] = 8'b11100000;
assign hamming[3721] = 8'b11100000;
assign hamming[3722] = 8'b11100001;
assign hamming[3723] = 8'b11100000;
assign hamming[3724] = 8'b11100001;
assign hamming[3725] = 8'b11100000;
assign hamming[3726] = 8'b11100001;
assign hamming[3727] = 8'b11100001;
assign hamming[3728] = 8'b11100010;
assign hamming[3729] = 8'b11100010;
assign hamming[3730] = 8'b11100010;
assign hamming[3731] = 8'b11100011;
assign hamming[3732] = 8'b11100010;
assign hamming[3733] = 8'b11100011;
assign hamming[3734] = 8'b11100011;
assign hamming[3735] = 8'b11100011;
assign hamming[3736] = 8'b11100010;
assign hamming[3737] = 8'b11100000;
assign hamming[3738] = 8'b11100110;
assign hamming[3739] = 8'b11101010;
assign hamming[3740] = 8'b11101011;
assign hamming[3741] = 8'b11100111;
assign hamming[3742] = 8'b11100001;
assign hamming[3743] = 8'b11100011;
assign hamming[3744] = 8'b11100101;
assign hamming[3745] = 8'b11100100;
assign hamming[3746] = 8'b11100100;
assign hamming[3747] = 8'b11100100;
assign hamming[3748] = 8'b11100101;
assign hamming[3749] = 8'b11100101;
assign hamming[3750] = 8'b11100101;
assign hamming[3751] = 8'b11100100;
assign hamming[3752] = 8'b11101100;
assign hamming[3753] = 8'b11100000;
assign hamming[3754] = 8'b11100110;
assign hamming[3755] = 8'b11100100;
assign hamming[3756] = 8'b11100101;
assign hamming[3757] = 8'b11100111;
assign hamming[3758] = 8'b11100001;
assign hamming[3759] = 8'b11101101;
assign hamming[3760] = 8'b11100010;
assign hamming[3761] = 8'b11101110;
assign hamming[3762] = 8'b11100110;
assign hamming[3763] = 8'b11100100;
assign hamming[3764] = 8'b11100101;
assign hamming[3765] = 8'b11100111;
assign hamming[3766] = 8'b11101111;
assign hamming[3767] = 8'b11100011;
assign hamming[3768] = 8'b11100110;
assign hamming[3769] = 8'b11100111;
assign hamming[3770] = 8'b11100110;
assign hamming[3771] = 8'b11100110;
assign hamming[3772] = 8'b11100111;
assign hamming[3773] = 8'b11100111;
assign hamming[3774] = 8'b11100110;
assign hamming[3775] = 8'b11100111;
assign hamming[3776] = 8'b11101000;
assign hamming[3777] = 8'b11101001;
assign hamming[3778] = 8'b11101000;
assign hamming[3779] = 8'b11101000;
assign hamming[3780] = 8'b11101001;
assign hamming[3781] = 8'b11101001;
assign hamming[3782] = 8'b11101000;
assign hamming[3783] = 8'b11101001;
assign hamming[3784] = 8'b11101100;
assign hamming[3785] = 8'b11100000;
assign hamming[3786] = 8'b11101000;
assign hamming[3787] = 8'b11101010;
assign hamming[3788] = 8'b11101011;
assign hamming[3789] = 8'b11101001;
assign hamming[3790] = 8'b11100001;
assign hamming[3791] = 8'b11101101;
assign hamming[3792] = 8'b11100010;
assign hamming[3793] = 8'b11101110;
assign hamming[3794] = 8'b11101000;
assign hamming[3795] = 8'b11101010;
assign hamming[3796] = 8'b11101011;
assign hamming[3797] = 8'b11101001;
assign hamming[3798] = 8'b11101111;
assign hamming[3799] = 8'b11100011;
assign hamming[3800] = 8'b11101011;
assign hamming[3801] = 8'b11101010;
assign hamming[3802] = 8'b11101010;
assign hamming[3803] = 8'b11101010;
assign hamming[3804] = 8'b11101011;
assign hamming[3805] = 8'b11101011;
assign hamming[3806] = 8'b11101011;
assign hamming[3807] = 8'b11101010;
assign hamming[3808] = 8'b11101100;
assign hamming[3809] = 8'b11101110;
assign hamming[3810] = 8'b11101000;
assign hamming[3811] = 8'b11100100;
assign hamming[3812] = 8'b11100101;
assign hamming[3813] = 8'b11101001;
assign hamming[3814] = 8'b11101111;
assign hamming[3815] = 8'b11101101;
assign hamming[3816] = 8'b11101100;
assign hamming[3817] = 8'b11101100;
assign hamming[3818] = 8'b11101100;
assign hamming[3819] = 8'b11101101;
assign hamming[3820] = 8'b11101100;
assign hamming[3821] = 8'b11101101;
assign hamming[3822] = 8'b11101101;
assign hamming[3823] = 8'b11101101;
assign hamming[3824] = 8'b11101110;
assign hamming[3825] = 8'b11101110;
assign hamming[3826] = 8'b11101111;
assign hamming[3827] = 8'b11101110;
assign hamming[3828] = 8'b11101111;
assign hamming[3829] = 8'b11101110;
assign hamming[3830] = 8'b11101111;
assign hamming[3831] = 8'b11101111;
assign hamming[3832] = 8'b11101100;
assign hamming[3833] = 8'b11101110;
assign hamming[3834] = 8'b11100110;
assign hamming[3835] = 8'b11101010;
assign hamming[3836] = 8'b11101011;
assign hamming[3837] = 8'b11100111;
assign hamming[3838] = 8'b11101111;
assign hamming[3839] = 8'b11101101;
assign hamming[3840] = 8'b11110000;
assign hamming[3841] = 8'b11110010;
assign hamming[3842] = 8'b11110100;
assign hamming[3843] = 8'b11111000;
assign hamming[3844] = 8'b11111001;
assign hamming[3845] = 8'b11110101;
assign hamming[3846] = 8'b11110011;
assign hamming[3847] = 8'b11110001;
assign hamming[3848] = 8'b11110000;
assign hamming[3849] = 8'b11110000;
assign hamming[3850] = 8'b11110000;
assign hamming[3851] = 8'b11110001;
assign hamming[3852] = 8'b11110000;
assign hamming[3853] = 8'b11110001;
assign hamming[3854] = 8'b11110001;
assign hamming[3855] = 8'b11110001;
assign hamming[3856] = 8'b11110010;
assign hamming[3857] = 8'b11110010;
assign hamming[3858] = 8'b11110011;
assign hamming[3859] = 8'b11110010;
assign hamming[3860] = 8'b11110011;
assign hamming[3861] = 8'b11110010;
assign hamming[3862] = 8'b11110011;
assign hamming[3863] = 8'b11110011;
assign hamming[3864] = 8'b11110000;
assign hamming[3865] = 8'b11110010;
assign hamming[3866] = 8'b11111010;
assign hamming[3867] = 8'b11110110;
assign hamming[3868] = 8'b11110111;
assign hamming[3869] = 8'b11111011;
assign hamming[3870] = 8'b11110011;
assign hamming[3871] = 8'b11110001;
assign hamming[3872] = 8'b11110100;
assign hamming[3873] = 8'b11110101;
assign hamming[3874] = 8'b11110100;
assign hamming[3875] = 8'b11110100;
assign hamming[3876] = 8'b11110101;
assign hamming[3877] = 8'b11110101;
assign hamming[3878] = 8'b11110100;
assign hamming[3879] = 8'b11110101;
assign hamming[3880] = 8'b11110000;
assign hamming[3881] = 8'b11111100;
assign hamming[3882] = 8'b11110100;
assign hamming[3883] = 8'b11110110;
assign hamming[3884] = 8'b11110111;
assign hamming[3885] = 8'b11110101;
assign hamming[3886] = 8'b11111101;
assign hamming[3887] = 8'b11110001;
assign hamming[3888] = 8'b11111110;
assign hamming[3889] = 8'b11110010;
assign hamming[3890] = 8'b11110100;
assign hamming[3891] = 8'b11110110;
assign hamming[3892] = 8'b11110111;
assign hamming[3893] = 8'b11110101;
assign hamming[3894] = 8'b11110011;
assign hamming[3895] = 8'b11111111;
assign hamming[3896] = 8'b11110111;
assign hamming[3897] = 8'b11110110;
assign hamming[3898] = 8'b11110110;
assign hamming[3899] = 8'b11110110;
assign hamming[3900] = 8'b11110111;
assign hamming[3901] = 8'b11110111;
assign hamming[3902] = 8'b11110111;
assign hamming[3903] = 8'b11110110;
assign hamming[3904] = 8'b11111001;
assign hamming[3905] = 8'b11111000;
assign hamming[3906] = 8'b11111000;
assign hamming[3907] = 8'b11111000;
assign hamming[3908] = 8'b11111001;
assign hamming[3909] = 8'b11111001;
assign hamming[3910] = 8'b11111001;
assign hamming[3911] = 8'b11111000;
assign hamming[3912] = 8'b11110000;
assign hamming[3913] = 8'b11111100;
assign hamming[3914] = 8'b11111010;
assign hamming[3915] = 8'b11111000;
assign hamming[3916] = 8'b11111001;
assign hamming[3917] = 8'b11111011;
assign hamming[3918] = 8'b11111101;
assign hamming[3919] = 8'b11110001;
assign hamming[3920] = 8'b11111110;
assign hamming[3921] = 8'b11110010;
assign hamming[3922] = 8'b11111010;
assign hamming[3923] = 8'b11111000;
assign hamming[3924] = 8'b11111001;
assign hamming[3925] = 8'b11111011;
assign hamming[3926] = 8'b11110011;
assign hamming[3927] = 8'b11111111;
assign hamming[3928] = 8'b11111010;
assign hamming[3929] = 8'b11111011;
assign hamming[3930] = 8'b11111010;
assign hamming[3931] = 8'b11111010;
assign hamming[3932] = 8'b11111011;
assign hamming[3933] = 8'b11111011;
assign hamming[3934] = 8'b11111010;
assign hamming[3935] = 8'b11111011;
assign hamming[3936] = 8'b11111110;
assign hamming[3937] = 8'b11111100;
assign hamming[3938] = 8'b11110100;
assign hamming[3939] = 8'b11111000;
assign hamming[3940] = 8'b11111001;
assign hamming[3941] = 8'b11110101;
assign hamming[3942] = 8'b11111101;
assign hamming[3943] = 8'b11111111;
assign hamming[3944] = 8'b11111100;
assign hamming[3945] = 8'b11111100;
assign hamming[3946] = 8'b11111101;
assign hamming[3947] = 8'b11111100;
assign hamming[3948] = 8'b11111101;
assign hamming[3949] = 8'b11111100;
assign hamming[3950] = 8'b11111101;
assign hamming[3951] = 8'b11111101;
assign hamming[3952] = 8'b11111110;
assign hamming[3953] = 8'b11111110;
assign hamming[3954] = 8'b11111110;
assign hamming[3955] = 8'b11111111;
assign hamming[3956] = 8'b11111110;
assign hamming[3957] = 8'b11111111;
assign hamming[3958] = 8'b11111111;
assign hamming[3959] = 8'b11111111;
assign hamming[3960] = 8'b11111110;
assign hamming[3961] = 8'b11111100;
assign hamming[3962] = 8'b11111010;
assign hamming[3963] = 8'b11110110;
assign hamming[3964] = 8'b11110111;
assign hamming[3965] = 8'b11111011;
assign hamming[3966] = 8'b11111101;
assign hamming[3967] = 8'b11111111;
assign hamming[3968] = 8'b01110000;
assign hamming[3969] = 8'b11111111;
assign hamming[3970] = 8'b11111111;
assign hamming[3971] = 8'b11111111;
assign hamming[3972] = 8'b11111111;
assign hamming[3973] = 8'b11111111;
assign hamming[3974] = 8'b11111111;
assign hamming[3975] = 8'b01110001;
assign hamming[3976] = 8'b11110000;
assign hamming[3977] = 8'b11100000;
assign hamming[3978] = 8'b11010000;
assign hamming[3979] = 8'b10110000;
assign hamming[3980] = 8'b10110001;
assign hamming[3981] = 8'b11010001;
assign hamming[3982] = 8'b11100001;
assign hamming[3983] = 8'b11110001;
assign hamming[3984] = 8'b11100010;
assign hamming[3985] = 8'b11110010;
assign hamming[3986] = 8'b10110010;
assign hamming[3987] = 8'b11010010;
assign hamming[3988] = 8'b11010011;
assign hamming[3989] = 8'b10110011;
assign hamming[3990] = 8'b11110011;
assign hamming[3991] = 8'b11100011;
assign hamming[3992] = 8'b11111111;
assign hamming[3993] = 8'b01110010;
assign hamming[3994] = 8'b11111111;
assign hamming[3995] = 8'b11111111;
assign hamming[3996] = 8'b11111111;
assign hamming[3997] = 8'b11111111;
assign hamming[3998] = 8'b01110011;
assign hamming[3999] = 8'b11111111;
assign hamming[4000] = 8'b11010100;
assign hamming[4001] = 8'b10110100;
assign hamming[4002] = 8'b11110100;
assign hamming[4003] = 8'b11100100;
assign hamming[4004] = 8'b11100101;
assign hamming[4005] = 8'b11110101;
assign hamming[4006] = 8'b10110101;
assign hamming[4007] = 8'b11010101;
assign hamming[4008] = 8'b11111111;
assign hamming[4009] = 8'b11111111;
assign hamming[4010] = 8'b01110100;
assign hamming[4011] = 8'b11111111;
assign hamming[4012] = 8'b11111111;
assign hamming[4013] = 8'b01110101;
assign hamming[4014] = 8'b11111111;
assign hamming[4015] = 8'b11111111;
assign hamming[4016] = 8'b11111111;
assign hamming[4017] = 8'b11111111;
assign hamming[4018] = 8'b11111111;
assign hamming[4019] = 8'b01110110;
assign hamming[4020] = 8'b01110111;
assign hamming[4021] = 8'b11111111;
assign hamming[4022] = 8'b11111111;
assign hamming[4023] = 8'b11111111;
assign hamming[4024] = 8'b10110110;
assign hamming[4025] = 8'b11010110;
assign hamming[4026] = 8'b11100110;
assign hamming[4027] = 8'b11110110;
assign hamming[4028] = 8'b11110111;
assign hamming[4029] = 8'b11100111;
assign hamming[4030] = 8'b11010111;
assign hamming[4031] = 8'b10110111;
assign hamming[4032] = 8'b10111000;
assign hamming[4033] = 8'b11011000;
assign hamming[4034] = 8'b11101000;
assign hamming[4035] = 8'b11111000;
assign hamming[4036] = 8'b11111001;
assign hamming[4037] = 8'b11101001;
assign hamming[4038] = 8'b11011001;
assign hamming[4039] = 8'b10111001;
assign hamming[4040] = 8'b11111111;
assign hamming[4041] = 8'b11111111;
assign hamming[4042] = 8'b11111111;
assign hamming[4043] = 8'b01111000;
assign hamming[4044] = 8'b01111001;
assign hamming[4045] = 8'b11111111;
assign hamming[4046] = 8'b11111111;
assign hamming[4047] = 8'b11111111;
assign hamming[4048] = 8'b11111111;
assign hamming[4049] = 8'b11111111;
assign hamming[4050] = 8'b01111010;
assign hamming[4051] = 8'b11111111;
assign hamming[4052] = 8'b11111111;
assign hamming[4053] = 8'b01111011;
assign hamming[4054] = 8'b11111111;
assign hamming[4055] = 8'b11111111;
assign hamming[4056] = 8'b11011010;
assign hamming[4057] = 8'b10111010;
assign hamming[4058] = 8'b11111010;
assign hamming[4059] = 8'b11101010;
assign hamming[4060] = 8'b11101011;
assign hamming[4061] = 8'b11111011;
assign hamming[4062] = 8'b10111011;
assign hamming[4063] = 8'b11011011;
assign hamming[4064] = 8'b11111111;
assign hamming[4065] = 8'b01111100;
assign hamming[4066] = 8'b11111111;
assign hamming[4067] = 8'b11111111;
assign hamming[4068] = 8'b11111111;
assign hamming[4069] = 8'b11111111;
assign hamming[4070] = 8'b01111101;
assign hamming[4071] = 8'b11111111;
assign hamming[4072] = 8'b11101100;
assign hamming[4073] = 8'b11111100;
assign hamming[4074] = 8'b10111100;
assign hamming[4075] = 8'b11011100;
assign hamming[4076] = 8'b11011101;
assign hamming[4077] = 8'b10111101;
assign hamming[4078] = 8'b11111101;
assign hamming[4079] = 8'b11101101;
assign hamming[4080] = 8'b11111110;
assign hamming[4081] = 8'b11101110;
assign hamming[4082] = 8'b11011110;
assign hamming[4083] = 8'b10111110;
assign hamming[4084] = 8'b10111111;
assign hamming[4085] = 8'b11011111;
assign hamming[4086] = 8'b11101111;
assign hamming[4087] = 8'b11111111;
assign hamming[4088] = 8'b01111110;
assign hamming[4089] = 8'b11111111;
assign hamming[4090] = 8'b11111111;
assign hamming[4091] = 8'b11111111;
assign hamming[4092] = 8'b11111111;
assign hamming[4093] = 8'b11111111;
assign hamming[4094] = 8'b11111111;
assign hamming[4095] = 8'b01111111;

input [11:0] datain;
output [7:0] dataout;

assign dataout = hamming[datain];

endmodule