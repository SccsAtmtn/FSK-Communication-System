module HammingCode(datain, dataout);

wire [11:0] hamming[255:0];
assign hamming[0] = 12'b000000000000;
assign hamming[1] = 12'b000000000111;
assign hamming[2] = 12'b000000011001;
assign hamming[3] = 12'b000000011110;
assign hamming[4] = 12'b000000101010;
assign hamming[5] = 12'b000000101101;
assign hamming[6] = 12'b000000110011;
assign hamming[7] = 12'b000000110100;
assign hamming[8] = 12'b000001001011;
assign hamming[9] = 12'b000001001100;
assign hamming[10] = 12'b000001010010;
assign hamming[11] = 12'b000001010101;
assign hamming[12] = 12'b000001100001;
assign hamming[13] = 12'b000001100110;
assign hamming[14] = 12'b000001111000;
assign hamming[15] = 12'b000001111111;
assign hamming[16] = 12'b000110000001;
assign hamming[17] = 12'b000110000110;
assign hamming[18] = 12'b000110011000;
assign hamming[19] = 12'b000110011111;
assign hamming[20] = 12'b000110101011;
assign hamming[21] = 12'b000110101100;
assign hamming[22] = 12'b000110110010;
assign hamming[23] = 12'b000110110101;
assign hamming[24] = 12'b000111001010;
assign hamming[25] = 12'b000111001101;
assign hamming[26] = 12'b000111010011;
assign hamming[27] = 12'b000111010100;
assign hamming[28] = 12'b000111100000;
assign hamming[29] = 12'b000111100111;
assign hamming[30] = 12'b000111111001;
assign hamming[31] = 12'b000111111110;
assign hamming[32] = 12'b001010000010;
assign hamming[33] = 12'b001010000101;
assign hamming[34] = 12'b001010011011;
assign hamming[35] = 12'b001010011100;
assign hamming[36] = 12'b001010101000;
assign hamming[37] = 12'b001010101111;
assign hamming[38] = 12'b001010110001;
assign hamming[39] = 12'b001010110110;
assign hamming[40] = 12'b001011001001;
assign hamming[41] = 12'b001011001110;
assign hamming[42] = 12'b001011010000;
assign hamming[43] = 12'b001011010111;
assign hamming[44] = 12'b001011100011;
assign hamming[45] = 12'b001011100100;
assign hamming[46] = 12'b001011111010;
assign hamming[47] = 12'b001011111101;
assign hamming[48] = 12'b001100000011;
assign hamming[49] = 12'b001100000100;
assign hamming[50] = 12'b001100011010;
assign hamming[51] = 12'b001100011101;
assign hamming[52] = 12'b001100101001;
assign hamming[53] = 12'b001100101110;
assign hamming[54] = 12'b001100110000;
assign hamming[55] = 12'b001100110111;
assign hamming[56] = 12'b001101001000;
assign hamming[57] = 12'b001101001111;
assign hamming[58] = 12'b001101010001;
assign hamming[59] = 12'b001101010110;
assign hamming[60] = 12'b001101100010;
assign hamming[61] = 12'b001101100101;
assign hamming[62] = 12'b001101111011;
assign hamming[63] = 12'b001101111100;
assign hamming[64] = 12'b010010000011;
assign hamming[65] = 12'b010010000100;
assign hamming[66] = 12'b010010011010;
assign hamming[67] = 12'b010010011101;
assign hamming[68] = 12'b010010101001;
assign hamming[69] = 12'b010010101110;
assign hamming[70] = 12'b010010110000;
assign hamming[71] = 12'b010010110111;
assign hamming[72] = 12'b010011001000;
assign hamming[73] = 12'b010011001111;
assign hamming[74] = 12'b010011010001;
assign hamming[75] = 12'b010011010110;
assign hamming[76] = 12'b010011100010;
assign hamming[77] = 12'b010011100101;
assign hamming[78] = 12'b010011111011;
assign hamming[79] = 12'b010011111100;
assign hamming[80] = 12'b010100000010;
assign hamming[81] = 12'b010100000101;
assign hamming[82] = 12'b010100011011;
assign hamming[83] = 12'b010100011100;
assign hamming[84] = 12'b010100101000;
assign hamming[85] = 12'b010100101111;
assign hamming[86] = 12'b010100110001;
assign hamming[87] = 12'b010100110110;
assign hamming[88] = 12'b010101001001;
assign hamming[89] = 12'b010101001110;
assign hamming[90] = 12'b010101010000;
assign hamming[91] = 12'b010101010111;
assign hamming[92] = 12'b010101100011;
assign hamming[93] = 12'b010101100100;
assign hamming[94] = 12'b010101111010;
assign hamming[95] = 12'b010101111101;
assign hamming[96] = 12'b011000000001;
assign hamming[97] = 12'b011000000110;
assign hamming[98] = 12'b011000011000;
assign hamming[99] = 12'b011000011111;
assign hamming[100] = 12'b011000101011;
assign hamming[101] = 12'b011000101100;
assign hamming[102] = 12'b011000110010;
assign hamming[103] = 12'b011000110101;
assign hamming[104] = 12'b011001001010;
assign hamming[105] = 12'b011001001101;
assign hamming[106] = 12'b011001010011;
assign hamming[107] = 12'b011001010100;
assign hamming[108] = 12'b011001100000;
assign hamming[109] = 12'b011001100111;
assign hamming[110] = 12'b011001111001;
assign hamming[111] = 12'b011001111110;
assign hamming[112] = 12'b011110000000;
assign hamming[113] = 12'b011110000111;
assign hamming[114] = 12'b011110011001;
assign hamming[115] = 12'b011110011110;
assign hamming[116] = 12'b011110101010;
assign hamming[117] = 12'b011110101101;
assign hamming[118] = 12'b011110110011;
assign hamming[119] = 12'b011110110100;
assign hamming[120] = 12'b011111001011;
assign hamming[121] = 12'b011111001100;
assign hamming[122] = 12'b011111010010;
assign hamming[123] = 12'b011111010101;
assign hamming[124] = 12'b011111100001;
assign hamming[125] = 12'b011111100110;
assign hamming[126] = 12'b011111111000;
assign hamming[127] = 12'b011111111111;
assign hamming[128] = 12'b100010001000;
assign hamming[129] = 12'b100010001111;
assign hamming[130] = 12'b100010010001;
assign hamming[131] = 12'b100010010110;
assign hamming[132] = 12'b100010100010;
assign hamming[133] = 12'b100010100101;
assign hamming[134] = 12'b100010111011;
assign hamming[135] = 12'b100010111100;
assign hamming[136] = 12'b100011000011;
assign hamming[137] = 12'b100011000100;
assign hamming[138] = 12'b100011011010;
assign hamming[139] = 12'b100011011101;
assign hamming[140] = 12'b100011101001;
assign hamming[141] = 12'b100011101110;
assign hamming[142] = 12'b100011110000;
assign hamming[143] = 12'b100011110111;
assign hamming[144] = 12'b100100001001;
assign hamming[145] = 12'b100100001110;
assign hamming[146] = 12'b100100010000;
assign hamming[147] = 12'b100100010111;
assign hamming[148] = 12'b100100100011;
assign hamming[149] = 12'b100100100100;
assign hamming[150] = 12'b100100111010;
assign hamming[151] = 12'b100100111101;
assign hamming[152] = 12'b100101000010;
assign hamming[153] = 12'b100101000101;
assign hamming[154] = 12'b100101011011;
assign hamming[155] = 12'b100101011100;
assign hamming[156] = 12'b100101101000;
assign hamming[157] = 12'b100101101111;
assign hamming[158] = 12'b100101110001;
assign hamming[159] = 12'b100101110110;
assign hamming[160] = 12'b101000001010;
assign hamming[161] = 12'b101000001101;
assign hamming[162] = 12'b101000010011;
assign hamming[163] = 12'b101000010100;
assign hamming[164] = 12'b101000100000;
assign hamming[165] = 12'b101000100111;
assign hamming[166] = 12'b101000111001;
assign hamming[167] = 12'b101000111110;
assign hamming[168] = 12'b101001000001;
assign hamming[169] = 12'b101001000110;
assign hamming[170] = 12'b101001011000;
assign hamming[171] = 12'b101001011111;
assign hamming[172] = 12'b101001101011;
assign hamming[173] = 12'b101001101100;
assign hamming[174] = 12'b101001110010;
assign hamming[175] = 12'b101001110101;
assign hamming[176] = 12'b101110001011;
assign hamming[177] = 12'b101110001100;
assign hamming[178] = 12'b101110010010;
assign hamming[179] = 12'b101110010101;
assign hamming[180] = 12'b101110100001;
assign hamming[181] = 12'b101110100110;
assign hamming[182] = 12'b101110111000;
assign hamming[183] = 12'b101110111111;
assign hamming[184] = 12'b101111000000;
assign hamming[185] = 12'b101111000111;
assign hamming[186] = 12'b101111011001;
assign hamming[187] = 12'b101111011110;
assign hamming[188] = 12'b101111101010;
assign hamming[189] = 12'b101111101101;
assign hamming[190] = 12'b101111110011;
assign hamming[191] = 12'b101111110100;
assign hamming[192] = 12'b110000001011;
assign hamming[193] = 12'b110000001100;
assign hamming[194] = 12'b110000010010;
assign hamming[195] = 12'b110000010101;
assign hamming[196] = 12'b110000100001;
assign hamming[197] = 12'b110000100110;
assign hamming[198] = 12'b110000111000;
assign hamming[199] = 12'b110000111111;
assign hamming[200] = 12'b110001000000;
assign hamming[201] = 12'b110001000111;
assign hamming[202] = 12'b110001011001;
assign hamming[203] = 12'b110001011110;
assign hamming[204] = 12'b110001101010;
assign hamming[205] = 12'b110001101101;
assign hamming[206] = 12'b110001110011;
assign hamming[207] = 12'b110001110100;
assign hamming[208] = 12'b110110001010;
assign hamming[209] = 12'b110110001101;
assign hamming[210] = 12'b110110010011;
assign hamming[211] = 12'b110110010100;
assign hamming[212] = 12'b110110100000;
assign hamming[213] = 12'b110110100111;
assign hamming[214] = 12'b110110111001;
assign hamming[215] = 12'b110110111110;
assign hamming[216] = 12'b110111000001;
assign hamming[217] = 12'b110111000110;
assign hamming[218] = 12'b110111011000;
assign hamming[219] = 12'b110111011111;
assign hamming[220] = 12'b110111101011;
assign hamming[221] = 12'b110111101100;
assign hamming[222] = 12'b110111110010;
assign hamming[223] = 12'b110111110101;
assign hamming[224] = 12'b111010001001;
assign hamming[225] = 12'b111010001110;
assign hamming[226] = 12'b111010010000;
assign hamming[227] = 12'b111010010111;
assign hamming[228] = 12'b111010100011;
assign hamming[229] = 12'b111010100100;
assign hamming[230] = 12'b111010111010;
assign hamming[231] = 12'b111010111101;
assign hamming[232] = 12'b111011000010;
assign hamming[233] = 12'b111011000101;
assign hamming[234] = 12'b111011011011;
assign hamming[235] = 12'b111011011100;
assign hamming[236] = 12'b111011101000;
assign hamming[237] = 12'b111011101111;
assign hamming[238] = 12'b111011110001;
assign hamming[239] = 12'b111011110110;
assign hamming[240] = 12'b111100001000;
assign hamming[241] = 12'b111100001111;
assign hamming[242] = 12'b111100010001;
assign hamming[243] = 12'b111100010110;
assign hamming[244] = 12'b111100100010;
assign hamming[245] = 12'b111100100101;
assign hamming[246] = 12'b111100111011;
assign hamming[247] = 12'b111100111100;
assign hamming[248] = 12'b111101000011;
assign hamming[249] = 12'b111101000100;
assign hamming[250] = 12'b111101011010;
assign hamming[251] = 12'b111101011101;
assign hamming[252] = 12'b111101101001;
assign hamming[253] = 12'b111101101110;
assign hamming[254] = 12'b111101110000;
assign hamming[255] = 12'b111101110111;

input [7:0] datain;
output [11:0] dataout;

assign dataout = hamming[datain];

endmodule